



//1014 * 36
//36 word length
//32 fraction length



module ln_ncpp_nvis_table(
    input [10-1:0] index, //0~1023
    output reg [36-1:0] table_out //36 word length, 32 fraction length
);

    always @(*) begin
        case (index)
            10'd0: table_out = 36'hddf95928a;
            10'd1: table_out = 36'hddfd4e0ac;
            10'd2: table_out = 36'hde0141f2b;
            10'd3: table_out = 36'hde0534e0e;
            10'd4: table_out = 36'hde0926d5c;
            10'd5: table_out = 36'hde0d17d1e;
            10'd6: table_out = 36'hde1107d5b;
            10'd7: table_out = 36'hde14f6e1b;
            10'd8: table_out = 36'hde18e4f65;
            10'd9: table_out = 36'hde1cd2140;
            10'd10: table_out = 36'hde20be3b6;
            10'd11: table_out = 36'hde24a96cc;
            10'd12: table_out = 36'hde2893a8b;
            10'd13: table_out = 36'hde2c7cefa;
            10'd14: table_out = 36'hde3065420;
            10'd15: table_out = 36'hde344ca05;
            10'd16: table_out = 36'hde38330b1;
            10'd17: table_out = 36'hde3c1882b;
            10'd18: table_out = 36'hde3ffd079;
            10'd19: table_out = 36'hde43e09a5;
            10'd20: table_out = 36'hde47c33b4;
            10'd21: table_out = 36'hde4ba4eae;
            10'd22: table_out = 36'hde4f85a9c;
            10'd23: table_out = 36'hde5365782;
            10'd24: table_out = 36'hde574456a;
            10'd25: table_out = 36'hde5b2245b;
            10'd26: table_out = 36'hde5eff45b;
            10'd27: table_out = 36'hde62db572;
            10'd28: table_out = 36'hde66b67a7;
            10'd29: table_out = 36'hde6a90b01;
            10'd30: table_out = 36'hde6e69f87;
            10'd31: table_out = 36'hde7242541;
            10'd32: table_out = 36'hde7619c35;
            10'd33: table_out = 36'hde79f046b;
            10'd34: table_out = 36'hde7dc5dea;
            10'd35: table_out = 36'hde819a8b8;
            10'd36: table_out = 36'hde856e4dd;
            10'd37: table_out = 36'hde8941260;
            10'd38: table_out = 36'hde8d13148;
            10'd39: table_out = 36'hde90e419c;
            10'd40: table_out = 36'hde94b4362;
            10'd41: table_out = 36'hde98836a2;
            10'd42: table_out = 36'hde9c51b62;
            10'd43: table_out = 36'hdea01f1aa;
            10'd44: table_out = 36'hdea3eb980;
            10'd45: table_out = 36'hdea7b72eb;
            10'd46: table_out = 36'hdeab81df2;
            10'd47: table_out = 36'hdeaf4ba9c;
            10'd48: table_out = 36'hdeb3148ef;
            10'd49: table_out = 36'hdeb6dc8f3;
            10'd50: table_out = 36'hdebaa3aae;
            10'd51: table_out = 36'hdebe69e27;
            10'd52: table_out = 36'hdec22f364;
            10'd53: table_out = 36'hdec5f3a6d;
            10'd54: table_out = 36'hdec9b7348;
            10'd55: table_out = 36'hdecd79dfb;
            10'd56: table_out = 36'hded13ba8e;
            10'd57: table_out = 36'hded4fc906;
            10'd58: table_out = 36'hded8bc96b;
            10'd59: table_out = 36'hdedc7bbc3;
            10'd60: table_out = 36'hdee03a015;
            10'd61: table_out = 36'hdee3f7667;
            10'd62: table_out = 36'hdee7b3ec0;
            10'd63: table_out = 36'hdeeb6f926;
            10'd64: table_out = 36'hdeef2a5a0;
            10'd65: table_out = 36'hdef2e4434;
            10'd66: table_out = 36'hdef69d4e9;
            10'd67: table_out = 36'hdefa557c5;
            10'd68: table_out = 36'hdefe0cccf;
            10'd69: table_out = 36'hdf01c340c;
            10'd70: table_out = 36'hdf0578d85;
            10'd71: table_out = 36'hdf092d93e;
            10'd72: table_out = 36'hdf0ce173e;
            10'd73: table_out = 36'hdf109478c;
            10'd74: table_out = 36'hdf1446a2d;
            10'd75: table_out = 36'hdf17f7f29;
            10'd76: table_out = 36'hdf1ba8686;
            10'd77: table_out = 36'hdf1f58049;
            10'd78: table_out = 36'hdf2306c79;
            10'd79: table_out = 36'hdf26b4b1c;
            10'd80: table_out = 36'hdf2a61c39;
            10'd81: table_out = 36'hdf2e0dfd5;
            10'd82: table_out = 36'hdf31b95f7;
            10'd83: table_out = 36'hdf3563ea6;
            10'd84: table_out = 36'hdf390d9e6;
            10'd85: table_out = 36'hdf3cb67bf;
            10'd86: table_out = 36'hdf405e837;
            10'd87: table_out = 36'hdf4405b52;
            10'd88: table_out = 36'hdf47ac119;
            10'd89: table_out = 36'hdf4b51991;
            10'd90: table_out = 36'hdf4ef64bf;
            10'd91: table_out = 36'hdf529a2aa;
            10'd92: table_out = 36'hdf563d358;
            10'd93: table_out = 36'hdf59df6cf;
            10'd94: table_out = 36'hdf5d80d15;
            10'd95: table_out = 36'hdf612162f;
            10'd96: table_out = 36'hdf64c1225;
            10'd97: table_out = 36'hdf68600fb;
            10'd98: table_out = 36'hdf6bfe2b8;
            10'd99: table_out = 36'hdf6f9b762;
            10'd100: table_out = 36'hdf7337efe;
            10'd101: table_out = 36'hdf76d3993;
            10'd102: table_out = 36'hdf7a6e726;
            10'd103: table_out = 36'hdf7e087bd;
            10'd104: table_out = 36'hdf81a1b5f;
            10'd105: table_out = 36'hdf853a210;
            10'd106: table_out = 36'hdf88d1bd7;
            10'd107: table_out = 36'hdf8c688b9;
            10'd108: table_out = 36'hdf8ffe8bc;
            10'd109: table_out = 36'hdf9393be6;
            10'd110: table_out = 36'hdf972823e;
            10'd111: table_out = 36'hdf9abbbc7;
            10'd112: table_out = 36'hdf9e4e889;
            10'd113: table_out = 36'hdfa1e0888;
            10'd114: table_out = 36'hdfa571bcc;
            10'd115: table_out = 36'hdfa902258;
            10'd116: table_out = 36'hdfac91c34;
            10'd117: table_out = 36'hdfb020963;
            10'd118: table_out = 36'hdfb3ae9ee;
            10'd119: table_out = 36'hdfb73bdd7;
            10'd120: table_out = 36'hdfbac8527;
            10'd121: table_out = 36'hdfbe53fe1;
            10'd122: table_out = 36'hdfc1dee0c;
            10'd123: table_out = 36'hdfc568fad;
            10'd124: table_out = 36'hdfc8f24c9;
            10'd125: table_out = 36'hdfcc7ad67;
            10'd126: table_out = 36'hdfd00298c;
            10'd127: table_out = 36'hdfd38993d;
            10'd128: table_out = 36'hdfd70fc7f;
            10'd129: table_out = 36'hdfda95358;
            10'd130: table_out = 36'hdfde19dcf;
            10'd131: table_out = 36'hdfe19dbe7;
            10'd132: table_out = 36'hdfe520da7;
            10'd133: table_out = 36'hdfe8a3313;
            10'd134: table_out = 36'hdfec24c32;
            10'd135: table_out = 36'hdfefa5909;
            10'd136: table_out = 36'hdff32599c;
            10'd137: table_out = 36'hdff6a4df2;
            10'd138: table_out = 36'hdffa23610;
            10'd139: table_out = 36'hdffda11fb;
            10'd140: table_out = 36'he0011e1b9;
            10'd141: table_out = 36'he0049a54e;
            10'd142: table_out = 36'he00815cc0;
            10'd143: table_out = 36'he00b90814;
            10'd144: table_out = 36'he00f0a750;
            10'd145: table_out = 36'he01283a79;
            10'd146: table_out = 36'he015fc194;
            10'd147: table_out = 36'he01973ca6;
            10'd148: table_out = 36'he01ceabb5;
            10'd149: table_out = 36'he02060ec5;
            10'd150: table_out = 36'he023d65dc;
            10'd151: table_out = 36'he0274b100;
            10'd152: table_out = 36'he02abf034;
            10'd153: table_out = 36'he02e3237f;
            10'd154: table_out = 36'he031a4ae5;
            10'd155: table_out = 36'he0351666c;
            10'd156: table_out = 36'he03887619;
            10'd157: table_out = 36'he03bf79f0;
            10'd158: table_out = 36'he03f671f7;
            10'd159: table_out = 36'he042d5e34;
            10'd160: table_out = 36'he04643eaa;
            10'd161: table_out = 36'he049b135f;
            10'd162: table_out = 36'he04d1dc59;
            10'd163: table_out = 36'he0508999b;
            10'd164: table_out = 36'he053f4b2c;
            10'd165: table_out = 36'he0575f110;
            10'd166: table_out = 36'he05ac8b4b;
            10'd167: table_out = 36'he05e319e4;
            10'd168: table_out = 36'he06199cdf;
            10'd169: table_out = 36'he06501441;
            10'd170: table_out = 36'he0686800f;
            10'd171: table_out = 36'he06bce04d;
            10'd172: table_out = 36'he06f33501;
            10'd173: table_out = 36'he07297e30;
            10'd174: table_out = 36'he075fbbde;
            10'd175: table_out = 36'he0795ee11;
            10'd176: table_out = 36'he07cc14cd;
            10'd177: table_out = 36'he08023017;
            10'd178: table_out = 36'he08383ff4;
            10'd179: table_out = 36'he086e4468;
            10'd180: table_out = 36'he08a43d79;
            10'd181: table_out = 36'he08da2b2c;
            10'd182: table_out = 36'he09100d84;
            10'd183: table_out = 36'he0945e487;
            10'd184: table_out = 36'he097bb03a;
            10'd185: table_out = 36'he09b170a2;
            10'd186: table_out = 36'he09e725c2;
            10'd187: table_out = 36'he0a1ccfa1;
            10'd188: table_out = 36'he0a526e42;
            10'd189: table_out = 36'he0a8801aa;
            10'd190: table_out = 36'he0abd89de;
            10'd191: table_out = 36'he0af306e3;
            10'd192: table_out = 36'he0b2878bd;
            10'd193: table_out = 36'he0b5ddf71;
            10'd194: table_out = 36'he0b933b04;
            10'd195: table_out = 36'he0bc88b7a;
            10'd196: table_out = 36'he0bfdd0d8;
            10'd197: table_out = 36'he0c330b23;
            10'd198: table_out = 36'he0c683a5f;
            10'd199: table_out = 36'he0c9d5e90;
            10'd200: table_out = 36'he0cd277bb;
            10'd201: table_out = 36'he0d0785e6;
            10'd202: table_out = 36'he0d3c8914;
            10'd203: table_out = 36'he0d71814a;
            10'd204: table_out = 36'he0da66e8c;
            10'd205: table_out = 36'he0ddb50df;
            10'd206: table_out = 36'he0e102848;
            10'd207: table_out = 36'he0e44f4cb;
            10'd208: table_out = 36'he0e79b66c;
            10'd209: table_out = 36'he0eae6d31;
            10'd210: table_out = 36'he0ee3191d;
            10'd211: table_out = 36'he0f17ba35;
            10'd212: table_out = 36'he0f4c507d;
            10'd213: table_out = 36'he0f80dbfa;
            10'd214: table_out = 36'he0fb55cb0;
            10'd215: table_out = 36'he0fe9d2a4;
            10'd216: table_out = 36'he101e3dda;
            10'd217: table_out = 36'he10529e56;
            10'd218: table_out = 36'he1086f41e;
            10'd219: table_out = 36'he10bb3f34;
            10'd220: table_out = 36'he10ef7f9e;
            10'd221: table_out = 36'he1123b561;
            10'd222: table_out = 36'he1157e07f;
            10'd223: table_out = 36'he118c00fe;
            10'd224: table_out = 36'he11c016e2;
            10'd225: table_out = 36'he11f4222f;
            10'd226: table_out = 36'he122822ea;
            10'd227: table_out = 36'he125c1916;
            10'd228: table_out = 36'he129004b9;
            10'd229: table_out = 36'he12c3e5d6;
            10'd230: table_out = 36'he12f7bc72;
            10'd231: table_out = 36'he132b8891;
            10'd232: table_out = 36'he135f4a36;
            10'd233: table_out = 36'he13930168;
            10'd234: table_out = 36'he13c6ae28;
            10'd235: table_out = 36'he13fa507d;
            10'd236: table_out = 36'he142de86a;
            10'd237: table_out = 36'he146175f3;
            10'd238: table_out = 36'he1494f91c;
            10'd239: table_out = 36'he14c871ea;
            10'd240: table_out = 36'he14fbe060;
            10'd241: table_out = 36'he152f4484;
            10'd242: table_out = 36'he15629e58;
            10'd243: table_out = 36'he1595ede2;
            10'd244: table_out = 36'he15c93325;
            10'd245: table_out = 36'he15fc6e25;
            10'd246: table_out = 36'he162f9ee7;
            10'd247: table_out = 36'he1662c56e;
            10'd248: table_out = 36'he1695e1bf;
            10'd249: table_out = 36'he16c8f3de;
            10'd250: table_out = 36'he16fbfbce;
            10'd251: table_out = 36'he172ef995;
            10'd252: table_out = 36'he1761ed35;
            10'd253: table_out = 36'he1794d6b3;
            10'd254: table_out = 36'he17c7b613;
            10'd255: table_out = 36'he17fa8b5a;
            10'd256: table_out = 36'he182d568a;
            10'd257: table_out = 36'he186017a8;
            10'd258: table_out = 36'he1892ceb8;
            10'd259: table_out = 36'he18c57bbe;
            10'd260: table_out = 36'he18f81ebe;
            10'd261: table_out = 36'he192ab7bc;
            10'd262: table_out = 36'he195d46bc;
            10'd263: table_out = 36'he198fcbc2;
            10'd264: table_out = 36'he19c246d1;
            10'd265: table_out = 36'he19f4b7ee;
            10'd266: table_out = 36'he1a271f1d;
            10'd267: table_out = 36'he1a597c61;
            10'd268: table_out = 36'he1a8bcfbf;
            10'd269: table_out = 36'he1abe1939;
            10'd270: table_out = 36'he1af058d5;
            10'd271: table_out = 36'he1b228e96;
            10'd272: table_out = 36'he1b54ba80;
            10'd273: table_out = 36'he1b86dc97;
            10'd274: table_out = 36'he1bb8f4de;
            10'd275: table_out = 36'he1beb0359;
            10'd276: table_out = 36'he1c1d080d;
            10'd277: table_out = 36'he1c4f02fd;
            10'd278: table_out = 36'he1c80f42d;
            10'd279: table_out = 36'he1cb2dba0;
            10'd280: table_out = 36'he1ce4b95b;
            10'd281: table_out = 36'he1d168d62;
            10'd282: table_out = 36'he1d4857b7;
            10'd283: table_out = 36'he1d7a185f;
            10'd284: table_out = 36'he1dabcf5d;
            10'd285: table_out = 36'he1ddd7cb6;
            10'd286: table_out = 36'he1e0f206d;
            10'd287: table_out = 36'he1e40ba86;
            10'd288: table_out = 36'he1e724b04;
            10'd289: table_out = 36'he1ea3d1ec;
            10'd290: table_out = 36'he1ed54f40;
            10'd291: table_out = 36'he1f06c305;
            10'd292: table_out = 36'he1f382d3f;
            10'd293: table_out = 36'he1f698df0;
            10'd294: table_out = 36'he1f9ae51d;
            10'd295: table_out = 36'he1fcc32c9;
            10'd296: table_out = 36'he1ffd76f9;
            10'd297: table_out = 36'he202eb1af;
            10'd298: table_out = 36'he205fe2ef;
            10'd299: table_out = 36'he20910abd;
            10'd300: table_out = 36'he20c2291d;
            10'd301: table_out = 36'he20f33e12;
            10'd302: table_out = 36'he212449a0;
            10'd303: table_out = 36'he21554bca;
            10'd304: table_out = 36'he21864494;
            10'd305: table_out = 36'he21b73402;
            10'd306: table_out = 36'he21e81a16;
            10'd307: table_out = 36'he2218f6d6;
            10'd308: table_out = 36'he2249ca44;
            10'd309: table_out = 36'he227a9463;
            10'd310: table_out = 36'he22ab5538;
            10'd311: table_out = 36'he22dc0cc6;
            10'd312: table_out = 36'he230cbb10;
            10'd313: table_out = 36'he233d601a;
            10'd314: table_out = 36'he236dfbe7;
            10'd315: table_out = 36'he239e8e7c;
            10'd316: table_out = 36'he23cf17db;
            10'd317: table_out = 36'he23ff9808;
            10'd318: table_out = 36'he24300f06;
            10'd319: table_out = 36'he24607cd9;
            10'd320: table_out = 36'he2490e185;
            10'd321: table_out = 36'he24c13d0c;
            10'd322: table_out = 36'he24f18f73;
            10'd323: table_out = 36'he2521d8bc;
            10'd324: table_out = 36'he255218ec;
            10'd325: table_out = 36'he25825005;
            10'd326: table_out = 36'he25b27e0b;
            10'd327: table_out = 36'he25e2a302;
            10'd328: table_out = 36'he2612beec;
            10'd329: table_out = 36'he2642d1ce;
            10'd330: table_out = 36'he2672dbaa;
            10'd331: table_out = 36'he26a2dc84;
            10'd332: table_out = 36'he26d2d45f;
            10'd333: table_out = 36'he2702c340;
            10'd334: table_out = 36'he2732a928;
            10'd335: table_out = 36'he2762861c;
            10'd336: table_out = 36'he27925a1f;
            10'd337: table_out = 36'he27c22533;
            10'd338: table_out = 36'he27f1e75e;
            10'd339: table_out = 36'he2821a0a1;
            10'd340: table_out = 36'he28515100;
            10'd341: table_out = 36'he2880f87e;
            10'd342: table_out = 36'he28b0971f;
            10'd343: table_out = 36'he28e02ce7;
            10'd344: table_out = 36'he290fb9d7;
            10'd345: table_out = 36'he293f3df4;
            10'd346: table_out = 36'he296eb941;
            10'd347: table_out = 36'he299e2bc2;
            10'd348: table_out = 36'he29cd9578;
            10'd349: table_out = 36'he29fcf668;
            10'd350: table_out = 36'he2a2c4e95;
            10'd351: table_out = 36'he2a5b9e02;
            10'd352: table_out = 36'he2a8ae4b3;
            10'd353: table_out = 36'he2aba22aa;
            10'd354: table_out = 36'he2ae957eb;
            10'd355: table_out = 36'he2b188479;
            10'd356: table_out = 36'he2b47a857;
            10'd357: table_out = 36'he2b76c389;
            10'd358: table_out = 36'he2ba5d611;
            10'd359: table_out = 36'he2bd4dff3;
            10'd360: table_out = 36'he2c03e131;
            10'd361: table_out = 36'he2c32d9d0;
            10'd362: table_out = 36'he2c61c9d3;
            10'd363: table_out = 36'he2c90b13b;
            10'd364: table_out = 36'he2cbf900e;
            10'd365: table_out = 36'he2cee664d;
            10'd366: table_out = 36'he2d1d33fc;
            10'd367: table_out = 36'he2d4bf91e;
            10'd368: table_out = 36'he2d7ab5b6;
            10'd369: table_out = 36'he2da969c7;
            10'd370: table_out = 36'he2dd81554;
            10'd371: table_out = 36'he2e06b862;
            10'd372: table_out = 36'he2e3552f1;
            10'd373: table_out = 36'he2e63e506;
            10'd374: table_out = 36'he2e926ea4;
            10'd375: table_out = 36'he2ec0efce;
            10'd376: table_out = 36'he2eef6887;
            10'd377: table_out = 36'he2f1dd8d1;
            10'd378: table_out = 36'he2f4c40b1;
            10'd379: table_out = 36'he2f7aa028;
            10'd380: table_out = 36'he2fa8f73b;
            10'd381: table_out = 36'he2fd745ec;
            10'd382: table_out = 36'he30058c3e;
            10'd383: table_out = 36'he3033ca34;
            10'd384: table_out = 36'he3061ffd1;
            10'd385: table_out = 36'he30902d18;
            10'd386: table_out = 36'he30be520d;
            10'd387: table_out = 36'he30ec6eb2;
            10'd388: table_out = 36'he311a830a;
            10'd389: table_out = 36'he31488f18;
            10'd390: table_out = 36'he317692df;
            10'd391: table_out = 36'he31a48e63;
            10'd392: table_out = 36'he31d281a5;
            10'd393: table_out = 36'he32006caa;
            10'd394: table_out = 36'he322e4f73;
            10'd395: table_out = 36'he325c2a05;
            10'd396: table_out = 36'he3289fc61;
            10'd397: table_out = 36'he32b7c68c;
            10'd398: table_out = 36'he32e58887;
            10'd399: table_out = 36'he33134256;
            10'd400: table_out = 36'he3340f3fb;
            10'd401: table_out = 36'he336e9d7a;
            10'd402: table_out = 36'he339c3ed5;
            10'd403: table_out = 36'he33c9d810;
            10'd404: table_out = 36'he33f7692d;
            10'd405: table_out = 36'he3424f22f;
            10'd406: table_out = 36'he34527318;
            10'd407: table_out = 36'he347febed;
            10'd408: table_out = 36'he34ad5cb0;
            10'd409: table_out = 36'he34dac563;
            10'd410: table_out = 36'he3508260a;
            10'd411: table_out = 36'he35357ea6;
            10'd412: table_out = 36'he3562cf3c;
            10'd413: table_out = 36'he359017ce;
            10'd414: table_out = 36'he35bd585f;
            10'd415: table_out = 36'he35ea90f2;
            10'd416: table_out = 36'he3617c189;
            10'd417: table_out = 36'he3644ea27;
            10'd418: table_out = 36'he36720acf;
            10'd419: table_out = 36'he369f2385;
            10'd420: table_out = 36'he36cc344a;
            10'd421: table_out = 36'he36f93d21;
            10'd422: table_out = 36'he37263e0e;
            10'd423: table_out = 36'he37533713;
            10'd424: table_out = 36'he37802832;
            10'd425: table_out = 36'he37ad1170;
            10'd426: table_out = 36'he37d9f2cd;
            10'd427: table_out = 36'he3806cc4e;
            10'd428: table_out = 36'he38339df5;
            10'd429: table_out = 36'he386067c4;
            10'd430: table_out = 36'he388d29bf;
            10'd431: table_out = 36'he38b9e3e7;
            10'd432: table_out = 36'he38e69641;
            10'd433: table_out = 36'he391340ce;
            10'd434: table_out = 36'he393fe392;
            10'd435: table_out = 36'he396c7e8e;
            10'd436: table_out = 36'he399911c6;
            10'd437: table_out = 36'he39c59d3d;
            10'd438: table_out = 36'he39f220f5;
            10'd439: table_out = 36'he3a1e9cf0;
            10'd440: table_out = 36'he3a4b1132;
            10'd441: table_out = 36'he3a777dbd;
            10'd442: table_out = 36'he3aa3e294;
            10'd443: table_out = 36'he3ad03fba;
            10'd444: table_out = 36'he3afc9531;
            10'd445: table_out = 36'he3b28e2fb;
            10'd446: table_out = 36'he3b55291c;
            10'd447: table_out = 36'he3b816796;
            10'd448: table_out = 36'he3bad9e6c;
            10'd449: table_out = 36'he3bd9cda1;
            10'd450: table_out = 36'he3c05f536;
            10'd451: table_out = 36'he3c32152f;
            10'd452: table_out = 36'he3c5e2d8f;
            10'd453: table_out = 36'he3c8a3e57;
            10'd454: table_out = 36'he3cb6478b;
            10'd455: table_out = 36'he3ce2492d;
            10'd456: table_out = 36'he3d0e4340;
            10'd457: table_out = 36'he3d3a35c6;
            10'd458: table_out = 36'he3d6620c2;
            10'd459: table_out = 36'he3d920436;
            10'd460: table_out = 36'he3dbde026;
            10'd461: table_out = 36'he3de9b493;
            10'd462: table_out = 36'he3e158181;
            10'd463: table_out = 36'he3e4146f1;
            10'd464: table_out = 36'he3e6d04e7;
            10'd465: table_out = 36'he3e98bb64;
            10'd466: table_out = 36'he3ec46a6c;
            10'd467: table_out = 36'he3ef01201;
            10'd468: table_out = 36'he3f1bb226;
            10'd469: table_out = 36'he3f474add;
            10'd470: table_out = 36'he3f72dc28;
            10'd471: table_out = 36'he3f9e660a;
            10'd472: table_out = 36'he3fc9e886;
            10'd473: table_out = 36'he3ff5639e;
            10'd474: table_out = 36'he4020d755;
            10'd475: table_out = 36'he404c43ad;
            10'd476: table_out = 36'he4077a8a9;
            10'd477: table_out = 36'he40a3064b;
            10'd478: table_out = 36'he40ce5c96;
            10'd479: table_out = 36'he40f9ab8b;
            10'd480: table_out = 36'he4124f32f;
            10'd481: table_out = 36'he41503382;
            10'd482: table_out = 36'he417b6c88;
            10'd483: table_out = 36'he41a69e43;
            10'd484: table_out = 36'he41d1c8b5;
            10'd485: table_out = 36'he41fcebe2;
            10'd486: table_out = 36'he422807ca;
            10'd487: table_out = 36'he42531c72;
            10'd488: table_out = 36'he427e29db;
            10'd489: table_out = 36'he42a93008;
            10'd490: table_out = 36'he42d42efa;
            10'd491: table_out = 36'he42ff26b6;
            10'd492: table_out = 36'he432a173c;
            10'd493: table_out = 36'he43550090;
            10'd494: table_out = 36'he437fe2b3;
            10'd495: table_out = 36'he43aabda9;
            10'd496: table_out = 36'he43d59173;
            10'd497: table_out = 36'he44005e15;
            10'd498: table_out = 36'he442b238f;
            10'd499: table_out = 36'he4455e1e6;
            10'd500: table_out = 36'he4480991b;
            10'd501: table_out = 36'he44ab4930;
            10'd502: table_out = 36'he44d5f228;
            10'd503: table_out = 36'he45009406;
            10'd504: table_out = 36'he452b2ecb;
            10'd505: table_out = 36'he4555c27a;
            10'd506: table_out = 36'he45804f16;
            10'd507: table_out = 36'he45aad4a0;
            10'd508: table_out = 36'he45d5531c;
            10'd509: table_out = 36'he45ffca8b;
            10'd510: table_out = 36'he462a3aef;
            10'd511: table_out = 36'he4654a44c;
            10'd512: table_out = 36'he467f06a3;
            10'd513: table_out = 36'he46a961f7;
            10'd514: table_out = 36'he46d3b64a;
            10'd515: table_out = 36'he46fe039f;
            10'd516: table_out = 36'he472849f7;
            10'd517: table_out = 36'he47528955;
            10'd518: table_out = 36'he477cc1bb;
            10'd519: table_out = 36'he47a6f32c;
            10'd520: table_out = 36'he47d11daa;
            10'd521: table_out = 36'he47fb4137;
            10'd522: table_out = 36'he48255dd5;
            10'd523: table_out = 36'he484f7387;
            10'd524: table_out = 36'he48798250;
            10'd525: table_out = 36'he48a38a30;
            10'd526: table_out = 36'he48cd8b2b;
            10'd527: table_out = 36'he48f78543;
            10'd528: table_out = 36'he4921787a;
            10'd529: table_out = 36'he494b64d2;
            10'd530: table_out = 36'he49754a4e;
            10'd531: table_out = 36'he499f28ef;
            10'd532: table_out = 36'he49c900b9;
            10'd533: table_out = 36'he49f2d1ad;
            10'd534: table_out = 36'he4a1c9bcd;
            10'd535: table_out = 36'he4a465f1d;
            10'd536: table_out = 36'he4a701b9d;
            10'd537: table_out = 36'he4a99d150;
            10'd538: table_out = 36'he4ac38039;
            10'd539: table_out = 36'he4aed2859;
            10'd540: table_out = 36'he4b16c9b3;
            10'd541: table_out = 36'he4b40644a;
            10'd542: table_out = 36'he4b69f81e;
            10'd543: table_out = 36'he4b938533;
            10'd544: table_out = 36'he4bbd0b8a;
            10'd545: table_out = 36'he4be68b27;
            10'd546: table_out = 36'he4c10040a;
            10'd547: table_out = 36'he4c397636;
            10'd548: table_out = 36'he4c62e1ae;
            10'd549: table_out = 36'he4c8c4673;
            10'd550: table_out = 36'he4cb5a488;
            10'd551: table_out = 36'he4cdefbee;
            10'd552: table_out = 36'he4d084ca9;
            10'd553: table_out = 36'he4d3196b9;
            10'd554: table_out = 36'he4d5ada22;
            10'd555: table_out = 36'he4d8416e6;
            10'd556: table_out = 36'he4dad4d06;
            10'd557: table_out = 36'he4dd67c84;
            10'd558: table_out = 36'he4dffa564;
            10'd559: table_out = 36'he4e28c7a6;
            10'd560: table_out = 36'he4e51e34d;
            10'd561: table_out = 36'he4e7af85c;
            10'd562: table_out = 36'he4ea406d4;
            10'd563: table_out = 36'he4ecd0eb7;
            10'd564: table_out = 36'he4ef61008;
            10'd565: table_out = 36'he4f1f0ac8;
            10'd566: table_out = 36'he4f47fefb;
            10'd567: table_out = 36'he4f70eca1;
            10'd568: table_out = 36'he4f99d3bd;
            10'd569: table_out = 36'he4fc2b451;
            10'd570: table_out = 36'he4feb8e5f;
            10'd571: table_out = 36'he501461e9;
            10'd572: table_out = 36'he503d2ef1;
            10'd573: table_out = 36'he5065f57a;
            10'd574: table_out = 36'he508eb585;
            10'd575: table_out = 36'he50b76f15;
            10'd576: table_out = 36'he50e0222b;
            10'd577: table_out = 36'he5108ceca;
            10'd578: table_out = 36'he513174f3;
            10'd579: table_out = 36'he515a14a9;
            10'd580: table_out = 36'he5182adee;
            10'd581: table_out = 36'he51ab40c3;
            10'd582: table_out = 36'he51d3cd2c;
            10'd583: table_out = 36'he51fc5329;
            10'd584: table_out = 36'he5224d2bd;
            10'd585: table_out = 36'he524d4bea;
            10'd586: table_out = 36'he5275beb2;
            10'd587: table_out = 36'he529e2b17;
            10'd588: table_out = 36'he52c6911a;
            10'd589: table_out = 36'he52eef0bf;
            10'd590: table_out = 36'he53174a07;
            10'd591: table_out = 36'he533f9cf3;
            10'd592: table_out = 36'he5367e987;
            10'd593: table_out = 36'he53902fc4;
            10'd594: table_out = 36'he53b86fab;
            10'd595: table_out = 36'he53e0a940;
            10'd596: table_out = 36'he5408dc83;
            10'd597: table_out = 36'he54310978;
            10'd598: table_out = 36'he5459301f;
            10'd599: table_out = 36'he5481507b;
            10'd600: table_out = 36'he54a96a8e;
            10'd601: table_out = 36'he54d17e5a;
            10'd602: table_out = 36'he54f98be1;
            10'd603: table_out = 36'he55219324;
            10'd604: table_out = 36'he55499427;
            10'd605: table_out = 36'he55718ee9;
            10'd606: table_out = 36'he5599836f;
            10'd607: table_out = 36'he55c171b9;
            10'd608: table_out = 36'he55e959c9;
            10'd609: table_out = 36'he56113ba2;
            10'd610: table_out = 36'he56391746;
            10'd611: table_out = 36'he5660ecb5;
            10'd612: table_out = 36'he5688bbf3;
            10'd613: table_out = 36'he56b08501;
            10'd614: table_out = 36'he56d847e1;
            10'd615: table_out = 36'he57000495;
            10'd616: table_out = 36'he5727bb1f;
            10'd617: table_out = 36'he574f6b81;
            10'd618: table_out = 36'he577715bd;
            10'd619: table_out = 36'he579eb9d4;
            10'd620: table_out = 36'he57c657c9;
            10'd621: table_out = 36'he57edef9d;
            10'd622: table_out = 36'he58158152;
            10'd623: table_out = 36'he583d0ceb;
            10'd624: table_out = 36'he58649269;
            10'd625: table_out = 36'he588c11ce;
            10'd626: table_out = 36'he58b38b1c;
            10'd627: table_out = 36'he58dafe54;
            10'd628: table_out = 36'he59026b79;
            10'd629: table_out = 36'he5929d28d;
            10'd630: table_out = 36'he59513391;
            10'd631: table_out = 36'he59788e87;
            10'd632: table_out = 36'he599fe371;
            10'd633: table_out = 36'he59c73252;
            10'd634: table_out = 36'he59ee7b2a;
            10'd635: table_out = 36'he5a15bdfb;
            10'd636: table_out = 36'he5a3cfac9;
            10'd637: table_out = 36'he5a643193;
            10'd638: table_out = 36'he5a8b625d;
            10'd639: table_out = 36'he5ab28d28;
            10'd640: table_out = 36'he5ad9b1f5;
            10'd641: table_out = 36'he5b00d0c8;
            10'd642: table_out = 36'he5b27e9a0;
            10'd643: table_out = 36'he5b4efc81;
            10'd644: table_out = 36'he5b76096d;
            10'd645: table_out = 36'he5b9d1064;
            10'd646: table_out = 36'he5bc41169;
            10'd647: table_out = 36'he5beb0c7d;
            10'd648: table_out = 36'he5c1201a3;
            10'd649: table_out = 36'he5c38f0dd;
            10'd650: table_out = 36'he5c5fda2b;
            10'd651: table_out = 36'he5c86bd90;
            10'd652: table_out = 36'he5cad9b0e;
            10'd653: table_out = 36'he5cd472a6;
            10'd654: table_out = 36'he5cfb445a;
            10'd655: table_out = 36'he5d22102c;
            10'd656: table_out = 36'he5d48d61e;
            10'd657: table_out = 36'he5d6f9631;
            10'd658: table_out = 36'he5d965068;
            10'd659: table_out = 36'he5dbd04c4;
            10'd660: table_out = 36'he5de3b346;
            10'd661: table_out = 36'he5e0a5bf2;
            10'd662: table_out = 36'he5e30fec7;
            10'd663: table_out = 36'he5e579bc9;
            10'd664: table_out = 36'he5e7e32f9;
            10'd665: table_out = 36'he5ea4c458;
            10'd666: table_out = 36'he5ecb4fe9;
            10'd667: table_out = 36'he5ef1d5ad;
            10'd668: table_out = 36'he5f1855a5;
            10'd669: table_out = 36'he5f3ecfd5;
            10'd670: table_out = 36'he5f65443c;
            10'd671: table_out = 36'he5f8bb2de;
            10'd672: table_out = 36'he5fb21bbc;
            10'd673: table_out = 36'he5fd87ed7;
            10'd674: table_out = 36'he5ffedc32;
            10'd675: table_out = 36'he602533cd;
            10'd676: table_out = 36'he604b85ab;
            10'd677: table_out = 36'he6071d1ce;
            10'd678: table_out = 36'he60981837;
            10'd679: table_out = 36'he60be58e8;
            10'd680: table_out = 36'he60e493e2;
            10'd681: table_out = 36'he610ac928;
            10'd682: table_out = 36'he6130f8ba;
            10'd683: table_out = 36'he6157229c;
            10'd684: table_out = 36'he617d46cd;
            10'd685: table_out = 36'he61a36551;
            10'd686: table_out = 36'he61c97e29;
            10'd687: table_out = 36'he61ef9156;
            10'd688: table_out = 36'he62159eda;
            10'd689: table_out = 36'he623ba6b7;
            10'd690: table_out = 36'he6261a8ee;
            10'd691: table_out = 36'he6287a582;
            10'd692: table_out = 36'he62ad9c74;
            10'd693: table_out = 36'he62d38dc5;
            10'd694: table_out = 36'he62f97977;
            10'd695: table_out = 36'he631f5f8c;
            10'd696: table_out = 36'he63454006;
            10'd697: table_out = 36'he636b1ae5;
            10'd698: table_out = 36'he6390f02d;
            10'd699: table_out = 36'he63b6bfde;
            10'd700: table_out = 36'he63dc89fa;
            10'd701: table_out = 36'he64024e83;
            10'd702: table_out = 36'he64280d7b;
            10'd703: table_out = 36'he644dc6e2;
            10'd704: table_out = 36'he64737abb;
            10'd705: table_out = 36'he64992908;
            10'd706: table_out = 36'he64bed1c9;
            10'd707: table_out = 36'he64e47501;
            10'd708: table_out = 36'he650a12b2;
            10'd709: table_out = 36'he652faadc;
            10'd710: table_out = 36'he65553d81;
            10'd711: table_out = 36'he657acaa4;
            10'd712: table_out = 36'he65a05245;
            10'd713: table_out = 36'he65c5d467;
            10'd714: table_out = 36'he65eb510b;
            10'd715: table_out = 36'he6610c832;
            10'd716: table_out = 36'he663639de;
            10'd717: table_out = 36'he665ba612;
            10'd718: table_out = 36'he66810ccd;
            10'd719: table_out = 36'he66a66e12;
            10'd720: table_out = 36'he66cbc9e3;
            10'd721: table_out = 36'he66f12041;
            10'd722: table_out = 36'he6716712e;
            10'd723: table_out = 36'he673bbcab;
            10'd724: table_out = 36'he676102ba;
            10'd725: table_out = 36'he6786435c;
            10'd726: table_out = 36'he67ab7e94;
            10'd727: table_out = 36'he67d0b462;
            10'd728: table_out = 36'he67f5e4c8;
            10'd729: table_out = 36'he681b0fc8;
            10'd730: table_out = 36'he68403563;
            10'd731: table_out = 36'he6865559c;
            10'd732: table_out = 36'he688a7072;
            10'd733: table_out = 36'he68af85e9;
            10'd734: table_out = 36'he68d49601;
            10'd735: table_out = 36'he68f9a0bd;
            10'd736: table_out = 36'he691ea61d;
            10'd737: table_out = 36'he6943a623;
            10'd738: table_out = 36'he6968a0d1;
            10'd739: table_out = 36'he698d9628;
            10'd740: table_out = 36'he69b2862a;
            10'd741: table_out = 36'he69d770d9;
            10'd742: table_out = 36'he69fc5635;
            10'd743: table_out = 36'he6a213641;
            10'd744: table_out = 36'he6a4610fe;
            10'd745: table_out = 36'he6a6ae66e;
            10'd746: table_out = 36'he6a8fb691;
            10'd747: table_out = 36'he6ab4816a;
            10'd748: table_out = 36'he6ad946fa;
            10'd749: table_out = 36'he6afe0743;
            10'd750: table_out = 36'he6b22c246;
            10'd751: table_out = 36'he6b477804;
            10'd752: table_out = 36'he6b6c2880;
            10'd753: table_out = 36'he6b90d3ba;
            10'd754: table_out = 36'he6bb579b5;
            10'd755: table_out = 36'he6bda1a71;
            10'd756: table_out = 36'he6bfeb5f0;
            10'd757: table_out = 36'he6c234c34;
            10'd758: table_out = 36'he6c47dd3e;
            10'd759: table_out = 36'he6c6c690f;
            10'd760: table_out = 36'he6c90efaa;
            10'd761: table_out = 36'he6cb5710f;
            10'd762: table_out = 36'he6cd9ed41;
            10'd763: table_out = 36'he6cfe6440;
            10'd764: table_out = 36'he6d22d60e;
            10'd765: table_out = 36'he6d4742ac;
            10'd766: table_out = 36'he6d6baa1d;
            10'd767: table_out = 36'he6d900c61;
            10'd768: table_out = 36'he6db4697a;
            10'd769: table_out = 36'he6dd8c169;
            10'd770: table_out = 36'he6dfd1431;
            10'd771: table_out = 36'he6e2161d1;
            10'd772: table_out = 36'he6e45aa4d;
            10'd773: table_out = 36'he6e69eda5;
            10'd774: table_out = 36'he6e8e2bda;
            10'd775: table_out = 36'he6eb264ef;
            10'd776: table_out = 36'he6ed698e4;
            10'd777: table_out = 36'he6efac7bb;
            10'd778: table_out = 36'he6f1ef176;
            10'd779: table_out = 36'he6f431616;
            10'd780: table_out = 36'he6f67359c;
            10'd781: table_out = 36'he6f8b500a;
            10'd782: table_out = 36'he6faf6561;
            10'd783: table_out = 36'he6fd375a3;
            10'd784: table_out = 36'he6ff780d2;
            10'd785: table_out = 36'he701b86ed;
            10'd786: table_out = 36'he703f87f8;
            10'd787: table_out = 36'he706383f3;
            10'd788: table_out = 36'he70877ae0;
            10'd789: table_out = 36'he70ab6cc0;
            10'd790: table_out = 36'he70cf5995;
            10'd791: table_out = 36'he70f34160;
            10'd792: table_out = 36'he71172423;
            10'd793: table_out = 36'he713b01de;
            10'd794: table_out = 36'he715eda94;
            10'd795: table_out = 36'he7182ae45;
            10'd796: table_out = 36'he71a67cf4;
            10'd797: table_out = 36'he71ca46a1;
            10'd798: table_out = 36'he71ee0b4e;
            10'd799: table_out = 36'he7211cafc;
            10'd800: table_out = 36'he723585ae;
            10'd801: table_out = 36'he72593b63;
            10'd802: table_out = 36'he727cec1e;
            10'd803: table_out = 36'he72a097df;
            10'd804: table_out = 36'he72c43ea9;
            10'd805: table_out = 36'he72e7e07d;
            10'd806: table_out = 36'he730b7d5b;
            10'd807: table_out = 36'he732f1546;
            10'd808: table_out = 36'he7352a83f;
            10'd809: table_out = 36'he73763647;
            10'd810: table_out = 36'he7399bf60;
            10'd811: table_out = 36'he73bd438a;
            10'd812: table_out = 36'he73e0c2c8;
            10'd813: table_out = 36'he74043d1a;
            10'd814: table_out = 36'he7427b283;
            10'd815: table_out = 36'he744b2302;
            10'd816: table_out = 36'he746e8e9b;
            10'd817: table_out = 36'he7491f54d;
            10'd818: table_out = 36'he74b5571b;
            10'd819: table_out = 36'he74d8b406;
            10'd820: table_out = 36'he74fc0c0f;
            10'd821: table_out = 36'he751f5f37;
            10'd822: table_out = 36'he7542ad80;
            10'd823: table_out = 36'he7565f6ec;
            10'd824: table_out = 36'he75893b7b;
            10'd825: table_out = 36'he75ac7b2e;
            10'd826: table_out = 36'he75cfb608;
            10'd827: table_out = 36'he75f2ec0a;
            10'd828: table_out = 36'he76161d34;
            10'd829: table_out = 36'he76394989;
            10'd830: table_out = 36'he765c7109;
            10'd831: table_out = 36'he767f93b5;
            10'd832: table_out = 36'he76a2b190;
            10'd833: table_out = 36'he76c5ca9b;
            10'd834: table_out = 36'he76e8ded6;
            10'd835: table_out = 36'he770bee44;
            10'd836: table_out = 36'he772ef8e4;
            10'd837: table_out = 36'he7751feba;
            10'd838: table_out = 36'he7774ffc6;
            10'd839: table_out = 36'he7797fc09;
            10'd840: table_out = 36'he77baf384;
            10'd841: table_out = 36'he77dde63a;
            10'd842: table_out = 36'he7800d42b;
            10'd843: table_out = 36'he7823bd59;
            10'd844: table_out = 36'he7846a1c4;
            10'd845: table_out = 36'he7869816f;
            10'd846: table_out = 36'he788c5c5a;
            10'd847: table_out = 36'he78af3286;
            10'd848: table_out = 36'he78d203f6;
            10'd849: table_out = 36'he78f4d0ab;
            10'd850: table_out = 36'he791798a4;
            10'd851: table_out = 36'he793a5be5;
            10'd852: table_out = 36'he795d1a6e;
            10'd853: table_out = 36'he797fd441;
            10'd854: table_out = 36'he79a2895e;
            10'd855: table_out = 36'he79c539c7;
            10'd856: table_out = 36'he79e7e57e;
            10'd857: table_out = 36'he7a0a8c83;
            10'd858: table_out = 36'he7a2d2ed8;
            10'd859: table_out = 36'he7a4fcc7e;
            10'd860: table_out = 36'he7a726576;
            10'd861: table_out = 36'he7a94f9c2;
            10'd862: table_out = 36'he7ab78963;
            10'd863: table_out = 36'he7ada145a;
            10'd864: table_out = 36'he7afc9aa9;
            10'd865: table_out = 36'he7b1f1c50;
            10'd866: table_out = 36'he7b419951;
            10'd867: table_out = 36'he7b6411ae;
            10'd868: table_out = 36'he7b868566;
            10'd869: table_out = 36'he7ba8f47d;
            10'd870: table_out = 36'he7bcb5ef2;
            10'd871: table_out = 36'he7bedc4c8;
            10'd872: table_out = 36'he7c1025ff;
            10'd873: table_out = 36'he7c328298;
            10'd874: table_out = 36'he7c54da96;
            10'd875: table_out = 36'he7c772df9;
            10'd876: table_out = 36'he7c997cc2;
            10'd877: table_out = 36'he7cbbc6f2;
            10'd878: table_out = 36'he7cde0c8c;
            10'd879: table_out = 36'he7d004d8f;
            10'd880: table_out = 36'he7d2289fe;
            10'd881: table_out = 36'he7d44c1d9;
            10'd882: table_out = 36'he7d66f522;
            10'd883: table_out = 36'he7d8923da;
            10'd884: table_out = 36'he7dab4e02;
            10'd885: table_out = 36'he7dcd739c;
            10'd886: table_out = 36'he7def94a8;
            10'd887: table_out = 36'he7e11b128;
            10'd888: table_out = 36'he7e33c91d;
            10'd889: table_out = 36'he7e55dc88;
            10'd890: table_out = 36'he7e77eb6a;
            10'd891: table_out = 36'he7e99f5c5;
            10'd892: table_out = 36'he7ebbfb9b;
            10'd893: table_out = 36'he7eddfceb;
            10'd894: table_out = 36'he7efff9b7;
            10'd895: table_out = 36'he7f21f201;
            10'd896: table_out = 36'he7f43e5c9;
            10'd897: table_out = 36'he7f65d512;
            10'd898: table_out = 36'he7f87bfdb;
            10'd899: table_out = 36'he7fa9a627;
            10'd900: table_out = 36'he7fcb87f6;
            10'd901: table_out = 36'he7fed6549;
            10'd902: table_out = 36'he800f3e23;
            10'd903: table_out = 36'he80311283;
            10'd904: table_out = 36'he8052e26b;
            10'd905: table_out = 36'he8074addd;
            10'd906: table_out = 36'he809674da;
            10'd907: table_out = 36'he80b83762;
            10'd908: table_out = 36'he80d9f576;
            10'd909: table_out = 36'he80fbaf19;
            10'd910: table_out = 36'he811d644b;
            10'd911: table_out = 36'he813f150e;
            10'd912: table_out = 36'he8160c162;
            10'd913: table_out = 36'he81826948;
            10'd914: table_out = 36'he81a40cc3;
            10'd915: table_out = 36'he81c5abd3;
            10'd916: table_out = 36'he81e74678;
            10'd917: table_out = 36'he8208dcb6;
            10'd918: table_out = 36'he822a6e8b;
            10'd919: table_out = 36'he824bfbfa;
            10'd920: table_out = 36'he826d8504;
            10'd921: table_out = 36'he828f09aa;
            10'd922: table_out = 36'he82b089ee;
            10'd923: table_out = 36'he82d205cf;
            10'd924: table_out = 36'he82f37d50;
            10'd925: table_out = 36'he8314f071;
            10'd926: table_out = 36'he83365f34;
            10'd927: table_out = 36'he8357c99a;
            10'd928: table_out = 36'he83792fa4;
            10'd929: table_out = 36'he839a9153;
            10'd930: table_out = 36'he83bbeea8;
            10'd931: table_out = 36'he83dd47a4;
            10'd932: table_out = 36'he83fe9c49;
            10'd933: table_out = 36'he841fec98;
            10'd934: table_out = 36'he84413892;
            10'd935: table_out = 36'he84628037;
            10'd936: table_out = 36'he8483c389;
            10'd937: table_out = 36'he84a5028a;
            10'd938: table_out = 36'he84c63d39;
            10'd939: table_out = 36'he84e77399;
            10'd940: table_out = 36'he8508a5ab;
            10'd941: table_out = 36'he8529d36f;
            10'd942: table_out = 36'he854afce7;
            10'd943: table_out = 36'he856c2214;
            10'd944: table_out = 36'he858d42f7;
            10'd945: table_out = 36'he85ae5f90;
            10'd946: table_out = 36'he85cf77e2;
            10'd947: table_out = 36'he85f08bee;
            10'd948: table_out = 36'he86119bb3;
            10'd949: table_out = 36'he8632a734;
            10'd950: table_out = 36'he8653ae72;
            10'd951: table_out = 36'he8674b16d;
            10'd952: table_out = 36'he8695b027;
            10'd953: table_out = 36'he86b6aaa1;
            10'd954: table_out = 36'he86d7a0dc;
            10'd955: table_out = 36'he86f892d9;
            10'd956: table_out = 36'he8719809a;
            10'd957: table_out = 36'he873a6a1e;
            10'd958: table_out = 36'he875b4f68;
            10'd959: table_out = 36'he877c3078;
            10'd960: table_out = 36'he879d0d50;
            10'd961: table_out = 36'he87bde5f0;
            10'd962: table_out = 36'he87deba5a;
            10'd963: table_out = 36'he87ff8a8f;
            10'd964: table_out = 36'he8820568f;
            10'd965: table_out = 36'he88411e5c;
            10'd966: table_out = 36'he8861e1f8;
            10'd967: table_out = 36'he8882a162;
            10'd968: table_out = 36'he88a35c9d;
            10'd969: table_out = 36'he88c413a9;
            10'd970: table_out = 36'he88e4c687;
            10'd971: table_out = 36'he89057538;
            10'd972: table_out = 36'he89261fbe;
            10'd973: table_out = 36'he8946c619;
            10'd974: table_out = 36'he8967684b;
            10'd975: table_out = 36'he89880654;
            10'd976: table_out = 36'he89a8a036;
            10'd977: table_out = 36'he89c935f2;
            10'd978: table_out = 36'he89e9c788;
            10'd979: table_out = 36'he8a0a54fa;
            10'd980: table_out = 36'he8a2ade49;
            10'd981: table_out = 36'he8a4b6376;
            10'd982: table_out = 36'he8a6be482;
            10'd983: table_out = 36'he8a8c616e;
            10'd984: table_out = 36'he8aacda3b;
            10'd985: table_out = 36'he8acd4eea;
            10'd986: table_out = 36'he8aedbf7c;
            10'd987: table_out = 36'he8b0e2bf3;
            10'd988: table_out = 36'he8b2e944e;
            10'd989: table_out = 36'he8b4ef890;
            10'd990: table_out = 36'he8b6f58b9;
            10'd991: table_out = 36'he8b8fb4cb;
            10'd992: table_out = 36'he8bb00cc6;
            10'd993: table_out = 36'he8bd060ab;
            10'd994: table_out = 36'he8bf0b07c;
            10'd995: table_out = 36'he8c10fc39;
            10'd996: table_out = 36'he8c3143e4;
            10'd997: table_out = 36'he8c51877d;
            10'd998: table_out = 36'he8c71c706;
            10'd999: table_out = 36'he8c92027f;
            10'd1000: table_out = 36'he8cb239ea;
            10'd1001: table_out = 36'he8cd26d47;
            10'd1002: table_out = 36'he8cf29c99;
            10'd1003: table_out = 36'he8d12c7de;
            10'd1004: table_out = 36'he8d32ef1a;
            10'd1005: table_out = 36'he8d53124c;
            10'd1006: table_out = 36'he8d733176;
            10'd1007: table_out = 36'he8d934c98;
            10'd1008: table_out = 36'he8db363b5;
            10'd1009: table_out = 36'he8dd376cc;
            10'd1010: table_out = 36'he8df385de;
            10'd1011: table_out = 36'he8e1390ee;
            10'd1012: table_out = 36'he8e3397fb;
            10'd1013: table_out = 36'he8e4fcaf1;
            default : table_out = 36'b0;
        endcase
    end



endmodule