


//1014 * 36
//36 word length
//32 fraction length



module ln_nvis_table(
    input [10-1:0] index, //0~1023
    output reg [36-1:0] table_out //36 word length, 32 fraction length
);

    always @(*) begin
        case (index)
            10'd0: table_out = 36'h94e12908f;
            10'd1: table_out = 36'h964e186e0;
            10'd2: table_out = 36'h979d249a7;
            10'd3: table_out = 36'h98d2d509f;
            10'd4: table_out = 36'h99f2bc03f;
            10'd5: table_out = 36'h9affb73dc;
            10'd6: table_out = 36'h9bfc1c7ee;
            10'd7: table_out = 36'h9ce9d9454;
            10'd8: table_out = 36'h9dca89b52;
            10'd9: table_out = 36'h9e9f898de;
            10'd10: table_out = 36'h9f6a00eba;
            10'd11: table_out = 36'ha02aee05f;
            10'd12: table_out = 36'ha0e32cbc6;
            10'd13: table_out = 36'ha1937c829;
            10'd14: table_out = 36'ha23c85128;
            10'd15: table_out = 36'ha2deda30b;
            10'd16: table_out = 36'ha37afeb84;
            10'd17: table_out = 36'ha41167171;
            10'd18: table_out = 36'ha4a27b59e;
            10'd19: table_out = 36'ha52e98de1;
            10'd20: table_out = 36'ha5b613bbe;
            10'd21: table_out = 36'ha63937f6d;
            10'd22: table_out = 36'ha6b84a7e2;
            10'd23: table_out = 36'ha7338a076;
            10'd24: table_out = 36'ha7ab2fc8b;
            10'd25: table_out = 36'ha81f7018a;
            10'd26: table_out = 36'ha8907af7e;
            10'd27: table_out = 36'ha8fe7c88c;
            10'd28: table_out = 36'ha9699d76a;
            10'd29: table_out = 36'ha9d20350b;
            10'd30: table_out = 36'haa37d0d8c;
            10'd31: table_out = 36'haa9b26494;
            10'd32: table_out = 36'haafc21924;
            10'd33: table_out = 36'hab5ade900;
            10'd34: table_out = 36'habb7773ad;
            10'd35: table_out = 36'hac1203d22;
            10'd36: table_out = 36'hac6a9b024;
            10'd37: table_out = 36'hacc152071;
            10'd38: table_out = 36'had163cca1;
            10'd39: table_out = 36'had696dfe3;
            10'd40: table_out = 36'hadbaf7385;
            10'd41: table_out = 36'hae0ae9060;
            10'd42: table_out = 36'hae5953010;
            10'd43: table_out = 36'haea643e26;
            10'd44: table_out = 36'haef1c9925;
            10'd45: table_out = 36'haf3bf137e;
            10'd46: table_out = 36'haf84c7465;
            10'd47: table_out = 36'hafcc5789d;
            10'd48: table_out = 36'hb012ad32f;
            10'd49: table_out = 36'hb057d2e15;
            10'd50: table_out = 36'hb09bd2ace;
            10'd51: table_out = 36'hb0deb62f2;
            10'd52: table_out = 36'hb120868b0;
            10'd53: table_out = 36'hb1614c747;
            10'd54: table_out = 36'hb1a110376;
            10'd55: table_out = 36'hb1dfd9be1;
            10'd56: table_out = 36'hb21db096f;
            10'd57: table_out = 36'hb25a9bfa2;
            10'd58: table_out = 36'hb296a2ce7;
            10'd59: table_out = 36'hb2d1cbae4;
            10'd60: table_out = 36'hb30c1ceba;
            10'd61: table_out = 36'hb3459c948;
            10'd62: table_out = 36'hb37e50767;
            10'd63: table_out = 36'hb3b63e222;
            10'd64: table_out = 36'hb3ed6aeeb;
            10'd65: table_out = 36'hb423dbfcd;
            10'd66: table_out = 36'hb45996396;
            10'd67: table_out = 36'hb48e9e605;
            10'd68: table_out = 36'hb4c2f8ff4;
            10'd69: table_out = 36'hb4f6aa777;
            10'd70: table_out = 36'hb529b7005;
            10'd71: table_out = 36'hb55c22a97;
            10'd72: table_out = 36'hb58df15c9;
            10'd73: table_out = 36'hb5bf26df1;
            10'd74: table_out = 36'hb5efc6d44;
            10'd75: table_out = 36'hb61fd4be5;
            10'd76: table_out = 36'hb64f54009;
            10'd77: table_out = 36'hb67e47e02;
            10'd78: table_out = 36'hb6acb385f;
            10'd79: table_out = 36'hb6da99ff9;
            10'd80: table_out = 36'hb707fe40b;
            10'd81: table_out = 36'hb734e3242;
            10'd82: table_out = 36'hb7614b6ce;
            10'd83: table_out = 36'hb78d39c73;
            10'd84: table_out = 36'hb7b8b0c9a;
            10'd85: table_out = 36'hb7e3b2f5c;
            10'd86: table_out = 36'hb80e42b93;
            10'd87: table_out = 36'hb838626e7;
            10'd88: table_out = 36'hb862145d7;
            10'd89: table_out = 36'hb88b5abca;
            10'd90: table_out = 36'hb8b437b18;
            10'd91: table_out = 36'hb8dcad511;
            10'd92: table_out = 36'hb904bda0f;
            10'd93: table_out = 36'hb92c6a979;
            10'd94: table_out = 36'hb953b61cf;
            10'd95: table_out = 36'hb97aa20b2;
            10'd96: table_out = 36'hb9a1302ee;
            10'd97: table_out = 36'hb9c76247f;
            10'd98: table_out = 36'hb9ed3a09c;
            10'd99: table_out = 36'hba12b91bd;
            10'd100: table_out = 36'hba37e11a0;
            10'd101: table_out = 36'hba5cb3951;
            10'd102: table_out = 36'hba8132133;
            10'd103: table_out = 36'hbaa55e101;
            10'd104: table_out = 36'hbac938fd8;
            10'd105: table_out = 36'hbaecc443b;
            10'd106: table_out = 36'hbb1001418;
            10'd107: table_out = 36'hbb32f14cc;
            10'd108: table_out = 36'hbb5595b2b;
            10'd109: table_out = 36'hbb77efb83;
            10'd110: table_out = 36'hbb9a0099f;
            10'd111: table_out = 36'hbbbbc98cc;
            10'd112: table_out = 36'hbbdd4bbe1;
            10'd113: table_out = 36'hbbfe8853c;
            10'd114: table_out = 36'hbc1f806cb;
            10'd115: table_out = 36'hbc403520e;
            10'd116: table_out = 36'hbc60a781b;
            10'd117: table_out = 36'hbc80d89a1;
            10'd118: table_out = 36'hbca0c96e9;
            10'd119: table_out = 36'hbcc07afdd;
            10'd120: table_out = 36'hbcdfee409;
            10'd121: table_out = 36'hbcff2429f;
            10'd122: table_out = 36'hbd1e1da75;
            10'd123: table_out = 36'hbd3cdba11;
            10'd124: table_out = 36'hbd5b5efa1;
            10'd125: table_out = 36'hbd79a8905;
            10'd126: table_out = 36'hbd97b93ce;
            10'd127: table_out = 36'hbdb591d42;
            10'd128: table_out = 36'hbdd33325c;
            10'd129: table_out = 36'hbdf09dfd0;
            10'd130: table_out = 36'hbe0dd320d;
            10'd131: table_out = 36'hbe2ad353d;
            10'd132: table_out = 36'hbe479f549;
            10'd133: table_out = 36'hbe6437ddb;
            10'd134: table_out = 36'hbe809da5e;
            10'd135: table_out = 36'hbe9cd1600;
            10'd136: table_out = 36'hbeb8d3bb6;
            10'd137: table_out = 36'hbed4a563b;
            10'd138: table_out = 36'hbef047011;
            10'd139: table_out = 36'hbf0bb9386;
            10'd140: table_out = 36'hbf26fcab3;
            10'd141: table_out = 36'hbf4211f7c;
            10'd142: table_out = 36'hbf5cf9b96;
            10'd143: table_out = 36'hbf77b4883;
            10'd144: table_out = 36'hbf9242f96;
            10'd145: table_out = 36'hbfaca59f4;
            10'd146: table_out = 36'hbfc6dd096;
            10'd147: table_out = 36'hbfe0e9c49;
            10'd148: table_out = 36'hbffacc5ad;
            10'd149: table_out = 36'hc0148553c;
            10'd150: table_out = 36'hc02e15344;
            10'd151: table_out = 36'hc0477c7ee;
            10'd152: table_out = 36'hc060bbb3c;
            10'd153: table_out = 36'hc079d3507;
            10'd154: table_out = 36'hc092c3d09;
            10'd155: table_out = 36'hc0ab8dad3;
            10'd156: table_out = 36'hc0c4315d6;
            10'd157: table_out = 36'hc0dcaf55f;
            10'd158: table_out = 36'hc0f50809c;
            10'd159: table_out = 36'hc10d3be98;
            10'd160: table_out = 36'hc1254b640;
            10'd161: table_out = 36'hc13d36e60;
            10'd162: table_out = 36'hc154feda8;
            10'd163: table_out = 36'hc16ca3aa9;
            10'd164: table_out = 36'hc18425bd7;
            10'd165: table_out = 36'hc19b8578a;
            10'd166: table_out = 36'hc1b2c33fe;
            10'd167: table_out = 36'hc1c9df755;
            10'd168: table_out = 36'hc1e0da796;
            10'd169: table_out = 36'hc1f7b4aae;
            10'd170: table_out = 36'hc20e6e670;
            10'd171: table_out = 36'hc22508098;
            10'd172: table_out = 36'hc23b81ec8;
            10'd173: table_out = 36'hc251dc68d;
            10'd174: table_out = 36'hc26817d5a;
            10'd175: table_out = 36'hc27e3488d;
            10'd176: table_out = 36'hc29432d6d;
            10'd177: table_out = 36'hc2aa1312d;
            10'd178: table_out = 36'hc2bfd58e9;
            10'd179: table_out = 36'hc2d57a9a9;
            10'd180: table_out = 36'hc2eb02860;
            10'd181: table_out = 36'hc3006d9ef;
            10'd182: table_out = 36'hc315bc321;
            10'd183: table_out = 36'hc32aee8af;
            10'd184: table_out = 36'hc34004f41;
            10'd185: table_out = 36'hc354ffb6a;
            10'd186: table_out = 36'hc369df1ad;
            10'd187: table_out = 36'hc37ea367a;
            10'd188: table_out = 36'hc3934ce31;
            10'd189: table_out = 36'hc3a7dbd21;
            10'd190: table_out = 36'hc3bc50788;
            10'd191: table_out = 36'hc3d0ab193;
            10'd192: table_out = 36'hc3e4ebf61;
            10'd193: table_out = 36'hc3f913500;
            10'd194: table_out = 36'hc40d21670;
            10'd195: table_out = 36'hc421167a1;
            10'd196: table_out = 36'hc434f2c75;
            10'd197: table_out = 36'hc448b68be;
            10'd198: table_out = 36'hc45c62042;
            10'd199: table_out = 36'hc46ff56b9;
            10'd200: table_out = 36'hc48370fcb;
            10'd201: table_out = 36'hc496d4f16;
            10'd202: table_out = 36'hc4aa21829;
            10'd203: table_out = 36'hc4bd56e86;
            10'd204: table_out = 36'hc4d0755a3;
            10'd205: table_out = 36'hc4e37d0eb;
            10'd206: table_out = 36'hc4f66e3ba;
            10'd207: table_out = 36'hc50949161;
            10'd208: table_out = 36'hc51c0dd28;
            10'd209: table_out = 36'hc52ebca48;
            10'd210: table_out = 36'hc54155bf0;
            10'd211: table_out = 36'hc553d9545;
            10'd212: table_out = 36'hc56647960;
            10'd213: table_out = 36'hc578a0b50;
            10'd214: table_out = 36'hc58ae4e18;
            10'd215: table_out = 36'hc59d144b3;
            10'd216: table_out = 36'hc5af2f210;
            10'd217: table_out = 36'hc5c135915;
            10'd218: table_out = 36'hc5d327c9e;
            10'd219: table_out = 36'hc5e505f7e;
            10'd220: table_out = 36'hc5f6d047e;
            10'd221: table_out = 36'hc60886e5d;
            10'd222: table_out = 36'hc61a29fd3;
            10'd223: table_out = 36'hc62bb9b8d;
            10'd224: table_out = 36'hc63d36431;
            10'd225: table_out = 36'hc64e9fc59;
            10'd226: table_out = 36'hc65ff669c;
            10'd227: table_out = 36'hc6713a583;
            10'd228: table_out = 36'hc6826bb93;
            10'd229: table_out = 36'hc6938ab46;
            10'd230: table_out = 36'hc6a497711;
            10'd231: table_out = 36'hc6b59215e;
            10'd232: table_out = 36'hc6c67ac91;
            10'd233: table_out = 36'hc6d751b07;
            10'd234: table_out = 36'hc6e816f15;
            10'd235: table_out = 36'hc6f8cab08;
            10'd236: table_out = 36'hc7096d127;
            10'd237: table_out = 36'hc719fe3b2;
            10'd238: table_out = 36'hc72a7e4df;
            10'd239: table_out = 36'hc73aed6e2;
            10'd240: table_out = 36'hc74b4bbe4;
            10'd241: table_out = 36'hc75b9960a;
            10'd242: table_out = 36'hc76bd6773;
            10'd243: table_out = 36'hc77c03234;
            10'd244: table_out = 36'hc78c1f85f;
            10'd245: table_out = 36'hc79c2bbff;
            10'd246: table_out = 36'hc7ac27f18;
            10'd247: table_out = 36'hc7bc143a9;
            10'd248: table_out = 36'hc7cbf0bab;
            10'd249: table_out = 36'hc7dbbd90f;
            10'd250: table_out = 36'hc7eb7adc5;
            10'd251: table_out = 36'hc7fb28bb2;
            10'd252: table_out = 36'hc80ac74b9;
            10'd253: table_out = 36'hc81a56ab5;
            10'd254: table_out = 36'hc829d6f7f;
            10'd255: table_out = 36'hc839484e7;
            10'd256: table_out = 36'hc848aacba;
            10'd257: table_out = 36'hc857fe8bf;
            10'd258: table_out = 36'hc86743ab8;
            10'd259: table_out = 36'hc8767a462;
            10'd260: table_out = 36'hc885a2776;
            10'd261: table_out = 36'hc894bc5a6;
            10'd262: table_out = 36'hc8a3c80a2;
            10'd263: table_out = 36'hc8b2c5a12;
            10'd264: table_out = 36'hc8c1b539c;
            10'd265: table_out = 36'hc8d096ee1;
            10'd266: table_out = 36'hc8df6ad7c;
            10'd267: table_out = 36'hc8ee31104;
            10'd268: table_out = 36'hc8fce9b0e;
            10'd269: table_out = 36'hc90b94d28;
            10'd270: table_out = 36'hc91a328dc;
            10'd271: table_out = 36'hc928c2fb1;
            10'd272: table_out = 36'hc93746329;
            10'd273: table_out = 36'hc945bc4c1;
            10'd274: table_out = 36'hc954255f5;
            10'd275: table_out = 36'hc96281839;
            10'd276: table_out = 36'hc970d0d01;
            10'd277: table_out = 36'hc97f135ba;
            10'd278: table_out = 36'hc98d493d0;
            10'd279: table_out = 36'hc99b728a7;
            10'd280: table_out = 36'hc9a98f5a5;
            10'd281: table_out = 36'hc9b79fc27;
            10'd282: table_out = 36'hc9c5a3d8b;
            10'd283: table_out = 36'hc9d39bb27;
            10'd284: table_out = 36'hc9e187650;
            10'd285: table_out = 36'hc9ef67059;
            10'd286: table_out = 36'hc9fd3aa8e;
            10'd287: table_out = 36'hca0b0263a;
            10'd288: table_out = 36'hca18be4a4;
            10'd289: table_out = 36'hca266e710;
            10'd290: table_out = 36'hca3412ebf;
            10'd291: table_out = 36'hca41abced;
            10'd292: table_out = 36'hca4f392d6;
            10'd293: table_out = 36'hca5cbb1b0;
            10'd294: table_out = 36'hca6a31aaf;
            10'd295: table_out = 36'hca779cf05;
            10'd296: table_out = 36'hca84fcfdf;
            10'd297: table_out = 36'hca9251e69;
            10'd298: table_out = 36'hca9f9bbcb;
            10'd299: table_out = 36'hcaacda929;
            10'd300: table_out = 36'hcaba0e7a8;
            10'd301: table_out = 36'hcac737865;
            10'd302: table_out = 36'hcad455c7e;
            10'd303: table_out = 36'hcae16950e;
            10'd304: table_out = 36'hcaee7232c;
            10'd305: table_out = 36'hcafb707ec;
            10'd306: table_out = 36'hcb0864461;
            10'd307: table_out = 36'hcb154d99b;
            10'd308: table_out = 36'hcb222c8a6;
            10'd309: table_out = 36'hcb2f0128e;
            10'd310: table_out = 36'hcb3bcb859;
            10'd311: table_out = 36'hcb488bb0e;
            10'd312: table_out = 36'hcb5541bb0;
            10'd313: table_out = 36'hcb61edb3f;
            10'd314: table_out = 36'hcb6e8faba;
            10'd315: table_out = 36'hcb7b27b1d;
            10'd316: table_out = 36'hcb87b5d62;
            10'd317: table_out = 36'hcb943a27f;
            10'd318: table_out = 36'hcba0b4b6b;
            10'd319: table_out = 36'hcbad25917;
            10'd320: table_out = 36'hcbb98cc75;
            10'd321: table_out = 36'hcbc5ea673;
            10'd322: table_out = 36'hcbd23e7fe;
            10'd323: table_out = 36'hcbde89200;
            10'd324: table_out = 36'hcbeaca560;
            10'd325: table_out = 36'hcbf702306;
            10'd326: table_out = 36'hcc0330bd4;
            10'd327: table_out = 36'hcc0f560ae;
            10'd328: table_out = 36'hcc1b72272;
            10'd329: table_out = 36'hcc27851ff;
            10'd330: table_out = 36'hcc338f031;
            10'd331: table_out = 36'hcc3f8fde2;
            10'd332: table_out = 36'hcc4b87bea;
            10'd333: table_out = 36'hcc5776b20;
            10'd334: table_out = 36'hcc635cc57;
            10'd335: table_out = 36'hcc6f3a063;
            10'd336: table_out = 36'hcc7b0e814;
            10'd337: table_out = 36'hcc86da43a;
            10'd338: table_out = 36'hcc929d5a1;
            10'd339: table_out = 36'hcc9e57d14;
            10'd340: table_out = 36'hccaa09b5e;
            10'd341: table_out = 36'hccb5b3147;
            10'd342: table_out = 36'hccc153f94;
            10'd343: table_out = 36'hccccec70a;
            10'd344: table_out = 36'hccd87c86c;
            10'd345: table_out = 36'hcce40447c;
            10'd346: table_out = 36'hccef83bf8;
            10'd347: table_out = 36'hccfafaf9f;
            10'd348: table_out = 36'hcd066a02e;
            10'd349: table_out = 36'hcd11d0e5f;
            10'd350: table_out = 36'hcd1d2faeb;
            10'd351: table_out = 36'hcd288668b;
            10'd352: table_out = 36'hcd33d51f4;
            10'd353: table_out = 36'hcd3f1bddb;
            10'd354: table_out = 36'hcd4a5aaf4;
            10'd355: table_out = 36'hcd55919f0;
            10'd356: table_out = 36'hcd60c0b7f;
            10'd357: table_out = 36'hcd6be8051;
            10'd358: table_out = 36'hcd7707912;
            10'd359: table_out = 36'hcd821f670;
            10'd360: table_out = 36'hcd8d2f913;
            10'd361: table_out = 36'hcd98381a7;
            10'd362: table_out = 36'hcda3390d2;
            10'd363: table_out = 36'hcdae3273b;
            10'd364: table_out = 36'hcdb924588;
            10'd365: table_out = 36'hcdc40ec5c;
            10'd366: table_out = 36'hcdcef1c59;
            10'd367: table_out = 36'hcdd9cd622;
            10'd368: table_out = 36'hcde4a1a56;
            10'd369: table_out = 36'hcdef6e994;
            10'd370: table_out = 36'hcdfa34479;
            10'd371: table_out = 36'hce04f2ba2;
            10'd372: table_out = 36'hce0fa9fa9;
            10'd373: table_out = 36'hce1a5a129;
            10'd374: table_out = 36'hce25030ba;
            10'd375: table_out = 36'hce2fa4ef3;
            10'd376: table_out = 36'hce3a3fc6b;
            10'd377: table_out = 36'hce44d39b7;
            10'd378: table_out = 36'hce4f6076b;
            10'd379: table_out = 36'hce59e6619;
            10'd380: table_out = 36'hce6465654;
            10'd381: table_out = 36'hce6edd8ab;
            10'd382: table_out = 36'hce794edaf;
            10'd383: table_out = 36'hce83b95ed;
            10'd384: table_out = 36'hce8e1d1f2;
            10'd385: table_out = 36'hce987a24c;
            10'd386: table_out = 36'hcea2d0785;
            10'd387: table_out = 36'hcead20227;
            10'd388: table_out = 36'hceb7692bc;
            10'd389: table_out = 36'hcec1ab9ca;
            10'd390: table_out = 36'hcecbe77da;
            10'd391: table_out = 36'hced61cd71;
            10'd392: table_out = 36'hcee04bb14;
            10'd393: table_out = 36'hceea74148;
            10'd394: table_out = 36'hcef49608e;
            10'd395: table_out = 36'hcefeb196a;
            10'd396: table_out = 36'hcf08c6c5c;
            10'd397: table_out = 36'hcf12d59e5;
            10'd398: table_out = 36'hcf1cde283;
            10'd399: table_out = 36'hcf26e06b5;
            10'd400: table_out = 36'hcf30dc6f8;
            10'd401: table_out = 36'hcf3ad23c9;
            10'd402: table_out = 36'hcf44c1da3;
            10'd403: table_out = 36'hcf4eab501;
            10'd404: table_out = 36'hcf588ea5d;
            10'd405: table_out = 36'hcf626be2e;
            10'd406: table_out = 36'hcf6c430ef;
            10'd407: table_out = 36'hcf7614314;
            10'd408: table_out = 36'hcf7fdf515;
            10'd409: table_out = 36'hcf89a4768;
            10'd410: table_out = 36'hcf9363a80;
            10'd411: table_out = 36'hcf9d1ced1;
            10'd412: table_out = 36'hcfa6d04cf;
            10'd413: table_out = 36'hcfb07dceb;
            10'd414: table_out = 36'hcfba25797;
            10'd415: table_out = 36'hcfc3c7544;
            10'd416: table_out = 36'hcfcd63660;
            10'd417: table_out = 36'hcfd6f9b5b;
            10'd418: table_out = 36'hcfe08a4a4;
            10'd419: table_out = 36'hcfea152a6;
            10'd420: table_out = 36'hcff39a5d0;
            10'd421: table_out = 36'hcffd19e8d;
            10'd422: table_out = 36'hd00693d48;
            10'd423: table_out = 36'hd0100826b;
            10'd424: table_out = 36'hd01976e60;
            10'd425: table_out = 36'hd022e0190;
            10'd426: table_out = 36'hd02c43c64;
            10'd427: table_out = 36'hd035a1f41;
            10'd428: table_out = 36'hd03efaa91;
            10'd429: table_out = 36'hd0484deb8;
            10'd430: table_out = 36'hd0519bc1b;
            10'd431: table_out = 36'hd05ae4320;
            10'd432: table_out = 36'hd0642742b;
            10'd433: table_out = 36'hd06d64f9e;
            10'd434: table_out = 36'hd0769d5dc;
            10'd435: table_out = 36'hd07fd0749;
            10'd436: table_out = 36'hd088fe443;
            10'd437: table_out = 36'hd09226d2e;
            10'd438: table_out = 36'hd09b4a267;
            10'd439: table_out = 36'hd0a468450;
            10'd440: table_out = 36'hd0ad81346;
            10'd441: table_out = 36'hd0b694fa8;
            10'd442: table_out = 36'hd0bfa39d3;
            10'd443: table_out = 36'hd0c8ad224;
            10'd444: table_out = 36'hd0d1b18f7;
            10'd445: table_out = 36'hd0dab0ea8;
            10'd446: table_out = 36'hd0e3ab392;
            10'd447: table_out = 36'hd0eca0810;
            10'd448: table_out = 36'hd0f590c7b;
            10'd449: table_out = 36'hd0fe7c12c;
            10'd450: table_out = 36'hd1076267d;
            10'd451: table_out = 36'hd11043cc5;
            10'd452: table_out = 36'hd1192045d;
            10'd453: table_out = 36'hd121f7d9a;
            10'd454: table_out = 36'hd12aca8d3;
            10'd455: table_out = 36'hd1339865f;
            10'd456: table_out = 36'hd13c61692;
            10'd457: table_out = 36'hd145259c1;
            10'd458: table_out = 36'hd14de5041;
            10'd459: table_out = 36'hd1569fa65;
            10'd460: table_out = 36'hd15f55880;
            10'd461: table_out = 36'hd16806ae5;
            10'd462: table_out = 36'hd170b31e6;
            10'd463: table_out = 36'hd1795add4;
            10'd464: table_out = 36'hd181fdf01;
            10'd465: table_out = 36'hd18a9c5bd;
            10'd466: table_out = 36'hd19336259;
            10'd467: table_out = 36'hd19bcb523;
            10'd468: table_out = 36'hd1a45be6a;
            10'd469: table_out = 36'hd1ace7e7e;
            10'd470: table_out = 36'hd1b56f5ad;
            10'd471: table_out = 36'hd1bdf2443;
            10'd472: table_out = 36'hd1c670a8e;
            10'd473: table_out = 36'hd1ceea8da;
            10'd474: table_out = 36'hd1d75ff74;
            10'd475: table_out = 36'hd1dfd0ea8;
            10'd476: table_out = 36'hd1e83d6c0;
            10'd477: table_out = 36'hd1f0a5807;
            10'd478: table_out = 36'hd1f9092c7;
            10'd479: table_out = 36'hd2016874b;
            10'd480: table_out = 36'hd209c35db;
            10'd481: table_out = 36'hd21219ec1;
            10'd482: table_out = 36'hd21a6c245;
            10'd483: table_out = 36'hd222ba0af;
            10'd484: table_out = 36'hd22b03a46;
            10'd485: table_out = 36'hd23348f53;
            10'd486: table_out = 36'hd23b8a01a;
            10'd487: table_out = 36'hd243c6ce4;
            10'd488: table_out = 36'hd24bff5f5;
            10'd489: table_out = 36'hd25433b93;
            10'd490: table_out = 36'hd25c63e03;
            10'd491: table_out = 36'hd2648fd8a;
            10'd492: table_out = 36'hd26cb7a6c;
            10'd493: table_out = 36'hd274db4ed;
            10'd494: table_out = 36'hd27cfad4f;
            10'd495: table_out = 36'hd285163d7;
            10'd496: table_out = 36'hd28d2d8c7;
            10'd497: table_out = 36'hd29540c61;
            10'd498: table_out = 36'hd29d4fee6;
            10'd499: table_out = 36'hd2a55b099;
            10'd500: table_out = 36'hd2ad621ba;
            10'd501: table_out = 36'hd2b56528a;
            10'd502: table_out = 36'hd2bd64349;
            10'd503: table_out = 36'hd2c55f437;
            10'd504: table_out = 36'hd2cd56594;
            10'd505: table_out = 36'hd2d54979f;
            10'd506: table_out = 36'hd2dd38a97;
            10'd507: table_out = 36'hd2e523eb9;
            10'd508: table_out = 36'hd2ed0b445;
            10'd509: table_out = 36'hd2f4eeb77;
            10'd510: table_out = 36'hd2fcce48e;
            10'd511: table_out = 36'hd304a9fc6;
            10'd512: table_out = 36'hd30c81d5c;
            10'd513: table_out = 36'hd31455d8c;
            10'd514: table_out = 36'hd31c26092;
            10'd515: table_out = 36'hd323f26aa;
            10'd516: table_out = 36'hd32bbb00f;
            10'd517: table_out = 36'hd3337fcfd;
            10'd518: table_out = 36'hd33b40dac;
            10'd519: table_out = 36'hd342fe259;
            10'd520: table_out = 36'hd34ab7b3d;
            10'd521: table_out = 36'hd3526d891;
            10'd522: table_out = 36'hd35a1fa8e;
            10'd523: table_out = 36'hd361ce16f;
            10'd524: table_out = 36'hd36978d6b;
            10'd525: table_out = 36'hd3711febb;
            10'd526: table_out = 36'hd378c3596;
            10'd527: table_out = 36'hd38063235;
            10'd528: table_out = 36'hd387ff4ce;
            10'd529: table_out = 36'hd38f97d9a;
            10'd530: table_out = 36'hd3972cccf;
            10'd531: table_out = 36'hd39ebe2a2;
            10'd532: table_out = 36'hd3a64bf4b;
            10'd533: table_out = 36'hd3add62ff;
            10'd534: table_out = 36'hd3b55cdf5;
            10'd535: table_out = 36'hd3bce0060;
            10'd536: table_out = 36'hd3c45fa76;
            10'd537: table_out = 36'hd3cbdbc6d;
            10'd538: table_out = 36'hd3d354677;
            10'd539: table_out = 36'hd3dac98ca;
            10'd540: table_out = 36'hd3e23b399;
            10'd541: table_out = 36'hd3e9a9718;
            10'd542: table_out = 36'hd3f11437a;
            10'd543: table_out = 36'hd3f87b8f2;
            10'd544: table_out = 36'hd3ffdf7b3;
            10'd545: table_out = 36'hd4073ffef;
            10'd546: table_out = 36'hd40e9d1d9;
            10'd547: table_out = 36'hd415f6da1;
            10'd548: table_out = 36'hd41d4d37b;
            10'd549: table_out = 36'hd424a0398;
            10'd550: table_out = 36'hd42befe27;
            10'd551: table_out = 36'hd4333c35c;
            10'd552: table_out = 36'hd43a85365;
            10'd553: table_out = 36'hd441cae73;
            10'd554: table_out = 36'hd4490d4b7;
            10'd555: table_out = 36'hd4504c660;
            10'd556: table_out = 36'hd4578839d;
            10'd557: table_out = 36'hd45ec0c9f;
            10'd558: table_out = 36'hd465f6194;
            10'd559: table_out = 36'hd46d282aa;
            10'd560: table_out = 36'hd47457011;
            10'd561: table_out = 36'hd47b829f7;
            10'd562: table_out = 36'hd482ab08a;
            10'd563: table_out = 36'hd489d03f8;
            10'd564: table_out = 36'hd490f246e;
            10'd565: table_out = 36'hd49811219;
            10'd566: table_out = 36'hd49f2cd28;
            10'd567: table_out = 36'hd4a6455c6;
            10'd568: table_out = 36'hd4ad5ac21;
            10'd569: table_out = 36'hd4b46d064;
            10'd570: table_out = 36'hd4bb7c2bd;
            10'd571: table_out = 36'hd4c288356;
            10'd572: table_out = 36'hd4c99125c;
            10'd573: table_out = 36'hd4d096ffb;
            10'd574: table_out = 36'hd4d799c5d;
            10'd575: table_out = 36'hd4de997ae;
            10'd576: table_out = 36'hd4e596218;
            10'd577: table_out = 36'hd4ec8fbc6;
            10'd578: table_out = 36'hd4f3864e3;
            10'd579: table_out = 36'hd4fa79d98;
            10'd580: table_out = 36'hd5016a610;
            10'd581: table_out = 36'hd50857e75;
            10'd582: table_out = 36'hd50f426f0;
            10'd583: table_out = 36'hd51629faa;
            10'd584: table_out = 36'hd51d0e8cd;
            10'd585: table_out = 36'hd523f0281;
            10'd586: table_out = 36'hd52acecf0;
            10'd587: table_out = 36'hd531aa841;
            10'd588: table_out = 36'hd5388349d;
            10'd589: table_out = 36'hd53f5922d;
            10'd590: table_out = 36'hd5462c118;
            10'd591: table_out = 36'hd54cfc185;
            10'd592: table_out = 36'hd553c939d;
            10'd593: table_out = 36'hd55a93786;
            10'd594: table_out = 36'hd5615ad69;
            10'd595: table_out = 36'hd5681f56b;
            10'd596: table_out = 36'hd56ee0fb3;
            10'd597: table_out = 36'hd5759fc69;
            10'd598: table_out = 36'hd57c5bbb2;
            10'd599: table_out = 36'hd58314db5;
            10'd600: table_out = 36'hd589cb297;
            10'd601: table_out = 36'hd5907ea7f;
            10'd602: table_out = 36'hd5972f591;
            10'd603: table_out = 36'hd59ddd3f4;
            10'd604: table_out = 36'hd5a4885cd;
            10'd605: table_out = 36'hd5ab30b40;
            10'd606: table_out = 36'hd5b1d6473;
            10'd607: table_out = 36'hd5b87918b;
            10'd608: table_out = 36'hd5bf192ab;
            10'd609: table_out = 36'hd5c5b67f8;
            10'd610: table_out = 36'hd5cc51197;
            10'd611: table_out = 36'hd5d2e8fab;
            10'd612: table_out = 36'hd5d97e259;
            10'd613: table_out = 36'hd5e0109c3;
            10'd614: table_out = 36'hd5e6a060e;
            10'd615: table_out = 36'hd5ed2d75c;
            10'd616: table_out = 36'hd5f3b7dd1;
            10'd617: table_out = 36'hd5fa3f990;
            10'd618: table_out = 36'hd600c4abc;
            10'd619: table_out = 36'hd60747176;
            10'd620: table_out = 36'hd60dc6de3;
            10'd621: table_out = 36'hd61444023;
            10'd622: table_out = 36'hd61abe85a;
            10'd623: table_out = 36'hd621366a9;
            10'd624: table_out = 36'hd627abb32;
            10'd625: table_out = 36'hd62e1e616;
            10'd626: table_out = 36'hd6348e778;
            10'd627: table_out = 36'hd63afbf78;
            10'd628: table_out = 36'hd64166e38;
            10'd629: table_out = 36'hd647cf3d9;
            10'd630: table_out = 36'hd64e3507b;
            10'd631: table_out = 36'hd65498440;
            10'd632: table_out = 36'hd65af8f48;
            10'd633: table_out = 36'hd661571b3;
            10'd634: table_out = 36'hd667b2ba1;
            10'd635: table_out = 36'hd66e0bd34;
            10'd636: table_out = 36'hd6746268a;
            10'd637: table_out = 36'hd67ab67c4;
            10'd638: table_out = 36'hd68108102;
            10'd639: table_out = 36'hd68757262;
            10'd640: table_out = 36'hd68da3c04;
            10'd641: table_out = 36'hd693ede08;
            10'd642: table_out = 36'hd69a3588c;
            10'd643: table_out = 36'hd6a07abb0;
            10'd644: table_out = 36'hd6a6bd792;
            10'd645: table_out = 36'hd6acfdc51;
            10'd646: table_out = 36'hd6b33ba0b;
            10'd647: table_out = 36'hd6b9770e0;
            10'd648: table_out = 36'hd6bfb00ed;
            10'd649: table_out = 36'hd6c5e6a50;
            10'd650: table_out = 36'hd6cc1ad27;
            10'd651: table_out = 36'hd6d24c990;
            10'd652: table_out = 36'hd6d87bfaa;
            10'd653: table_out = 36'hd6dea8f90;
            10'd654: table_out = 36'hd6e4d3962;
            10'd655: table_out = 36'hd6eafbd3c;
            10'd656: table_out = 36'hd6f121b3b;
            10'd657: table_out = 36'hd6f74537c;
            10'd658: table_out = 36'hd6fd6661d;
            10'd659: table_out = 36'hd7038533a;
            10'd660: table_out = 36'hd709a1aef;
            10'd661: table_out = 36'hd70fbbd5a;
            10'd662: table_out = 36'hd715d3a97;
            10'd663: table_out = 36'hd71be92c2;
            10'd664: table_out = 36'hd721fc5f6;
            10'd665: table_out = 36'hd7280d451;
            10'd666: table_out = 36'hd72e1bdee;
            10'd667: table_out = 36'hd734282e9;
            10'd668: table_out = 36'hd73a3235d;
            10'd669: table_out = 36'hd74039f66;
            10'd670: table_out = 36'hd7463f720;
            10'd671: table_out = 36'hd74c42aa5;
            10'd672: table_out = 36'hd75243a12;
            10'd673: table_out = 36'hd75842580;
            10'd674: table_out = 36'hd75e3ed0b;
            10'd675: table_out = 36'hd764390cd;
            10'd676: table_out = 36'hd76a310e2;
            10'd677: table_out = 36'hd77026d65;
            10'd678: table_out = 36'hd7761a66e;
            10'd679: table_out = 36'hd77c0bc19;
            10'd680: table_out = 36'hd781fae80;
            10'd681: table_out = 36'hd787e7dbe;
            10'd682: table_out = 36'hd78dd29eb;
            10'd683: table_out = 36'hd793bb323;
            10'd684: table_out = 36'hd799a197e;
            10'd685: table_out = 36'hd79f85d17;
            10'd686: table_out = 36'hd7a567e07;
            10'd687: table_out = 36'hd7ab47c67;
            10'd688: table_out = 36'hd7b125851;
            10'd689: table_out = 36'hd7b7011df;
            10'd690: table_out = 36'hd7bcda928;
            10'd691: table_out = 36'hd7c2b1e47;
            10'd692: table_out = 36'hd7c887154;
            10'd693: table_out = 36'hd7ce5a268;
            10'd694: table_out = 36'hd7d42b19b;
            10'd695: table_out = 36'hd7d9f9f07;
            10'd696: table_out = 36'hd7dfc6ac3;
            10'd697: table_out = 36'hd7e5914e8;
            10'd698: table_out = 36'hd7eb59d8f;
            10'd699: table_out = 36'hd7f1204d0;
            10'd700: table_out = 36'hd7f6e4ac2;
            10'd701: table_out = 36'hd7fca6f7d;
            10'd702: table_out = 36'hd8026731b;
            10'd703: table_out = 36'hd808255b1;
            10'd704: table_out = 36'hd80de1758;
            10'd705: table_out = 36'hd8139b828;
            10'd706: table_out = 36'hd81953838;
            10'd707: table_out = 36'hd81f097a0;
            10'd708: table_out = 36'hd824bd675;
            10'd709: table_out = 36'hd82a6f4d1;
            10'd710: table_out = 36'hd8301f2ca;
            10'd711: table_out = 36'hd835cd077;
            10'd712: table_out = 36'hd83b78dee;
            10'd713: table_out = 36'hd84122b47;
            10'd714: table_out = 36'hd846ca899;
            10'd715: table_out = 36'hd84c705f9;
            10'd716: table_out = 36'hd8521437f;
            10'd717: table_out = 36'hd857b6140;
            10'd718: table_out = 36'hd85d55f54;
            10'd719: table_out = 36'hd862f3dd0;
            10'd720: table_out = 36'hd8688fccb;
            10'd721: table_out = 36'hd86e29c5b;
            10'd722: table_out = 36'hd873c1c95;
            10'd723: table_out = 36'hd87957d90;
            10'd724: table_out = 36'hd87eebf61;
            10'd725: table_out = 36'hd8847e21e;
            10'd726: table_out = 36'hd88a0e5dd;
            10'd727: table_out = 36'hd88f9cab2;
            10'd728: table_out = 36'hd895290b5;
            10'd729: table_out = 36'hd89ab37f9;
            10'd730: table_out = 36'hd8a03c095;
            10'd731: table_out = 36'hd8a5c2a9c;
            10'd732: table_out = 36'hd8ab47626;
            10'd733: table_out = 36'hd8b0ca346;
            10'd734: table_out = 36'hd8b64b211;
            10'd735: table_out = 36'hd8bbca29c;
            10'd736: table_out = 36'hd8c1474fd;
            10'd737: table_out = 36'hd8c6c2947;
            10'd738: table_out = 36'hd8cc3bf8f;
            10'd739: table_out = 36'hd8d1b37ea;
            10'd740: table_out = 36'hd8d72926c;
            10'd741: table_out = 36'hd8dc9cf2a;
            10'd742: table_out = 36'hd8e20ee37;
            10'd743: table_out = 36'hd8e77efa9;
            10'd744: table_out = 36'hd8eced392;
            10'd745: table_out = 36'hd8f259a08;
            10'd746: table_out = 36'hd8f7c431e;
            10'd747: table_out = 36'hd8fd2cee7;
            10'd748: table_out = 36'hd90293d78;
            10'd749: table_out = 36'hd907f8ee5;
            10'd750: table_out = 36'hd90d5c340;
            10'd751: table_out = 36'hd912bda9e;
            10'd752: table_out = 36'hd9181d512;
            10'd753: table_out = 36'hd91d7b2b0;
            10'd754: table_out = 36'hd922d738a;
            10'd755: table_out = 36'hd928317b4;
            10'd756: table_out = 36'hd92d89f41;
            10'd757: table_out = 36'hd932e0a45;
            10'd758: table_out = 36'hd938358d2;
            10'd759: table_out = 36'hd93d88afb;
            10'd760: table_out = 36'hd942da0d3;
            10'd761: table_out = 36'hd94829a6d;
            10'd762: table_out = 36'hd94d777db;
            10'd763: table_out = 36'hd952c3931;
            10'd764: table_out = 36'hd9580de80;
            10'd765: table_out = 36'hd95d567dc;
            10'd766: table_out = 36'hd9629d557;
            10'd767: table_out = 36'hd967e2703;
            10'd768: table_out = 36'hd96d25cf2;
            10'd769: table_out = 36'hd97267737;
            10'd770: table_out = 36'hd977a75e4;
            10'd771: table_out = 36'hd97ce590b;
            10'd772: table_out = 36'hd982220bd;
            10'd773: table_out = 36'hd9875cd0e;
            10'd774: table_out = 36'hd98c95e0e;
            10'd775: table_out = 36'hd991cd3d0;
            10'd776: table_out = 36'hd99702e65;
            10'd777: table_out = 36'hd99c36ddf;
            10'd778: table_out = 36'hd9a16924f;
            10'd779: table_out = 36'hd9a699bc8;
            10'd780: table_out = 36'hd9abc8a5a;
            10'd781: table_out = 36'hd9b0f5e17;
            10'd782: table_out = 36'hd9b621711;
            10'd783: table_out = 36'hd9bb4b558;
            10'd784: table_out = 36'hd9c0738fe;
            10'd785: table_out = 36'hd9c59a214;
            10'd786: table_out = 36'hd9cabf0ab;
            10'd787: table_out = 36'hd9cfe24d4;
            10'd788: table_out = 36'hd9d503ea0;
            10'd789: table_out = 36'hd9da23e20;
            10'd790: table_out = 36'hd9df42364;
            10'd791: table_out = 36'hd9e45ee7f;
            10'd792: table_out = 36'hd9e979f7f;
            10'd793: table_out = 36'hd9ee93676;
            10'd794: table_out = 36'hd9f3ab374;
            10'd795: table_out = 36'hd9f8c168b;
            10'd796: table_out = 36'hd9fdd5fca;
            10'd797: table_out = 36'hda02e8f41;
            10'd798: table_out = 36'hda07fa502;
            10'd799: table_out = 36'hda0d0a11c;
            10'd800: table_out = 36'hda121839f;
            10'd801: table_out = 36'hda1724c9d;
            10'd802: table_out = 36'hda1c2fc24;
            10'd803: table_out = 36'hda2139245;
            10'd804: table_out = 36'hda2640f0f;
            10'd805: table_out = 36'hda2b47294;
            10'd806: table_out = 36'hda304bce1;
            10'd807: table_out = 36'hda354ee09;
            10'd808: table_out = 36'hda3a50619;
            10'd809: table_out = 36'hda3f50522;
            10'd810: table_out = 36'hda444eb34;
            10'd811: table_out = 36'hda494b85e;
            10'd812: table_out = 36'hda4e46caf;
            10'd813: table_out = 36'hda5340837;
            10'd814: table_out = 36'hda5838b05;
            10'd815: table_out = 36'hda5d2f529;
            10'd816: table_out = 36'hda62246b2;
            10'd817: table_out = 36'hda6717faf;
            10'd818: table_out = 36'hda6c0a02f;
            10'd819: table_out = 36'hda70fa842;
            10'd820: table_out = 36'hda75e97f7;
            10'd821: table_out = 36'hda7ad6f5c;
            10'd822: table_out = 36'hda7fc2e80;
            10'd823: table_out = 36'hda84ad573;
            10'd824: table_out = 36'hda8996443;
            10'd825: table_out = 36'hda8e7daff;
            10'd826: table_out = 36'hda93639b6;
            10'd827: table_out = 36'hda9848077;
            10'd828: table_out = 36'hda9d2af50;
            10'd829: table_out = 36'hdaa20c64f;
            10'd830: table_out = 36'hdaa6ec583;
            10'd831: table_out = 36'hdaabcacfc;
            10'd832: table_out = 36'hdab0a7cc6;
            10'd833: table_out = 36'hdab5834f1;
            10'd834: table_out = 36'hdaba5d58b;
            10'd835: table_out = 36'hdabf35ea2;
            10'd836: table_out = 36'hdac40d044;
            10'd837: table_out = 36'hdac8e2a80;
            10'd838: table_out = 36'hdacdb6d63;
            10'd839: table_out = 36'hdad2898fc;
            10'd840: table_out = 36'hdad75ad59;
            10'd841: table_out = 36'hdadc2aa88;
            10'd842: table_out = 36'hdae0f9096;
            10'd843: table_out = 36'hdae5c5f92;
            10'd844: table_out = 36'hdaea91789;
            10'd845: table_out = 36'hdaef5b889;
            10'd846: table_out = 36'hdaf4242a0;
            10'd847: table_out = 36'hdaf8eb5dc;
            10'd848: table_out = 36'hdafdb124a;
            10'd849: table_out = 36'hdb02757f7;
            10'd850: table_out = 36'hdb07386f2;
            10'd851: table_out = 36'hdb0bf9f48;
            10'd852: table_out = 36'hdb10ba106;
            10'd853: table_out = 36'hdb1578c3a;
            10'd854: table_out = 36'hdb1a360f0;
            10'd855: table_out = 36'hdb1ef1f38;
            10'd856: table_out = 36'hdb23ac71c;
            10'd857: table_out = 36'hdb28658ab;
            10'd858: table_out = 36'hdb2d1d3f3;
            10'd859: table_out = 36'hdb31d38ff;
            10'd860: table_out = 36'hdb36887de;
            10'd861: table_out = 36'hdb3b3c09c;
            10'd862: table_out = 36'hdb3fee346;
            10'd863: table_out = 36'hdb449efe9;
            10'd864: table_out = 36'hdb494e692;
            10'd865: table_out = 36'hdb4dfc74e;
            10'd866: table_out = 36'hdb52a922a;
            10'd867: table_out = 36'hdb5754732;
            10'd868: table_out = 36'hdb5bfe673;
            10'd869: table_out = 36'hdb60a6ffb;
            10'd870: table_out = 36'hdb654e3d4;
            10'd871: table_out = 36'hdb69f420d;
            10'd872: table_out = 36'hdb6e98ab2;
            10'd873: table_out = 36'hdb733bdcf;
            10'd874: table_out = 36'hdb77ddb70;
            10'd875: table_out = 36'hdb7c7e3a2;
            10'd876: table_out = 36'hdb811d672;
            10'd877: table_out = 36'hdb85bb3ec;
            10'd878: table_out = 36'hdb8a57c1c;
            10'd879: table_out = 36'hdb8ef2f0e;
            10'd880: table_out = 36'hdb938ccce;
            10'd881: table_out = 36'hdb982556a;
            10'd882: table_out = 36'hdb9cbc8ec;
            10'd883: table_out = 36'hdba152761;
            10'd884: table_out = 36'hdba5e70d6;
            10'd885: table_out = 36'hdbaa7a555;
            10'd886: table_out = 36'hdbaf0c4eb;
            10'd887: table_out = 36'hdbb39cfa4;
            10'd888: table_out = 36'hdbb82c58c;
            10'd889: table_out = 36'hdbbcba6af;
            10'd890: table_out = 36'hdbc147318;
            10'd891: table_out = 36'hdbc5d2ad3;
            10'd892: table_out = 36'hdbca5cded;
            10'd893: table_out = 36'hdbcee5c70;
            10'd894: table_out = 36'hdbd36d668;
            10'd895: table_out = 36'hdbd7f3be2;
            10'd896: table_out = 36'hdbdc78ce8;
            10'd897: table_out = 36'hdbe0fc986;
            10'd898: table_out = 36'hdbe57f1c7;
            10'd899: table_out = 36'hdbea005b8;
            10'd900: table_out = 36'hdbee80563;
            10'd901: table_out = 36'hdbf2ff0d4;
            10'd902: table_out = 36'hdbf77c816;
            10'd903: table_out = 36'hdbfbf8b35;
            10'd904: table_out = 36'hdc0073a3c;
            10'd905: table_out = 36'hdc04ed536;
            10'd906: table_out = 36'hdc0965c2e;
            10'd907: table_out = 36'hdc0ddcf2f;
            10'd908: table_out = 36'hdc1252e45;
            10'd909: table_out = 36'hdc16c797b;
            10'd910: table_out = 36'hdc1b3b0db;
            10'd911: table_out = 36'hdc1fad471;
            10'd912: table_out = 36'hdc241e448;
            10'd913: table_out = 36'hdc288e06a;
            10'd914: table_out = 36'hdc2cfc8e3;
            10'd915: table_out = 36'hdc3169dbe;
            10'd916: table_out = 36'hdc35d5f05;
            10'd917: table_out = 36'hdc3a40cc3;
            10'd918: table_out = 36'hdc3eaa703;
            10'd919: table_out = 36'hdc4312dcf;
            10'd920: table_out = 36'hdc477a133;
            10'd921: table_out = 36'hdc4be0139;
            10'd922: table_out = 36'hdc5044dec;
            10'd923: table_out = 36'hdc54a8755;
            10'd924: table_out = 36'hdc590ad81;
            10'd925: table_out = 36'hdc5d6c079;
            10'd926: table_out = 36'hdc61cc048;
            10'd927: table_out = 36'hdc662acf8;
            10'd928: table_out = 36'hdc6a88694;
            10'd929: table_out = 36'hdc6ee4d26;
            10'd930: table_out = 36'hdc73400b9;
            10'd931: table_out = 36'hdc779a157;
            10'd932: table_out = 36'hdc7bf2f09;
            10'd933: table_out = 36'hdc804a9dc;
            10'd934: table_out = 36'hdc84a11d7;
            10'd935: table_out = 36'hdc88f6707;
            10'd936: table_out = 36'hdc8d4a975;
            10'd937: table_out = 36'hdc919d92b;
            10'd938: table_out = 36'hdc95ef633;
            10'd939: table_out = 36'hdc9a40098;
            10'd940: table_out = 36'hdc9e8f863;
            10'd941: table_out = 36'hdca2ddd9e;
            10'd942: table_out = 36'hdca72b054;
            10'd943: table_out = 36'hdcab7708e;
            10'd944: table_out = 36'hdcafc1e57;
            10'd945: table_out = 36'hdcb40b9b7;
            10'd946: table_out = 36'hdcb8542ba;
            10'd947: table_out = 36'hdcbc9b969;
            10'd948: table_out = 36'hdcc0e1dcd;
            10'd949: table_out = 36'hdcc526ff0;
            10'd950: table_out = 36'hdcc96afdd;
            10'd951: table_out = 36'hdccdadd9c;
            10'd952: table_out = 36'hdcd1ef938;
            10'd953: table_out = 36'hdcd6302ba;
            10'd954: table_out = 36'hdcda6fa2c;
            10'd955: table_out = 36'hdcdeadf97;
            10'd956: table_out = 36'hdce2eb305;
            10'd957: table_out = 36'hdce727480;
            10'd958: table_out = 36'hdceb62410;
            10'd959: table_out = 36'hdcef9c1bf;
            10'd960: table_out = 36'hdcf3d4d98;
            10'd961: table_out = 36'hdcf80c7a3;
            10'd962: table_out = 36'hdcfc42fe9;
            10'd963: table_out = 36'hdd0078674;
            10'd964: table_out = 36'hdd04acb4d;
            10'd965: table_out = 36'hdd08dfe7e;
            10'd966: table_out = 36'hdd0d12010;
            10'd967: table_out = 36'hdd114300c;
            10'd968: table_out = 36'hdd1572e7b;
            10'd969: table_out = 36'hdd19a1b66;
            10'd970: table_out = 36'hdd1dcf6d7;
            10'd971: table_out = 36'hdd21fc0d7;
            10'd972: table_out = 36'hdd262796e;
            10'd973: table_out = 36'hdd2a520a6;
            10'd974: table_out = 36'hdd2e7b688;
            10'd975: table_out = 36'hdd32a3b1d;
            10'd976: table_out = 36'hdd36cae6e;
            10'd977: table_out = 36'hdd3af1083;
            10'd978: table_out = 36'hdd3f16167;
            10'd979: table_out = 36'hdd433a121;
            10'd980: table_out = 36'hdd475cfba;
            10'd981: table_out = 36'hdd4b7ed3c;
            10'd982: table_out = 36'hdd4f9f9af;
            10'd983: table_out = 36'hdd53bf51c;
            10'd984: table_out = 36'hdd57ddf8c;
            10'd985: table_out = 36'hdd5bfb907;
            10'd986: table_out = 36'hdd6018196;
            10'd987: table_out = 36'hdd6433942;
            10'd988: table_out = 36'hdd684e014;
            10'd989: table_out = 36'hdd6c67614;
            10'd990: table_out = 36'hdd707fb4b;
            10'd991: table_out = 36'hdd7496fc1;
            10'd992: table_out = 36'hdd78ad37f;
            10'd993: table_out = 36'hdd7cc268e;
            10'd994: table_out = 36'hdd80d68f5;
            10'd995: table_out = 36'hdd84e9abe;
            10'd996: table_out = 36'hdd88fbbf1;
            10'd997: table_out = 36'hdd8d0cc96;
            10'd998: table_out = 36'hdd911ccb6;
            10'd999: table_out = 36'hdd952bc59;
            10'd1000: table_out = 36'hdd9939b87;
            10'd1001: table_out = 36'hdd9d46a4a;
            10'd1002: table_out = 36'hdda1528a8;
            10'd1003: table_out = 36'hdda55d6ab;
            10'd1004: table_out = 36'hdda96745a;
            10'd1005: table_out = 36'hddad701bf;
            10'd1006: table_out = 36'hddb177ee0;
            10'd1007: table_out = 36'hddb57ebc7;
            10'd1008: table_out = 36'hddb98487b;
            10'd1009: table_out = 36'hddbd89505;
            10'd1010: table_out = 36'hddc18d16d;
            10'd1011: table_out = 36'hddc58fdba;
            10'd1012: table_out = 36'hddc9919f5;
            10'd1013: table_out = 36'hddcd185d1;
            default: table_out = 36'b0;
        endcase
    end


endmodule