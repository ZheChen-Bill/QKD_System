

//1229 * 36
//36 word length
//32 fraction length


module log2_1_p_table(
    input [11-1:0] index, //0~2047
    output reg [36-1:0] table_out //36 word length, 32 fraction length
);

    always @(*) begin
        case (index)
            11'd0: table_out = 36'head799f13;
            11'd1: table_out = 36'head3fe0e9;
            11'd2: table_out = 36'head0619b7;
            11'd3: table_out = 36'heaccc4979;
            11'd4: table_out = 36'heac92702d;
            11'd5: table_out = 36'heac588dd0;
            11'd6: table_out = 36'heac1ea25f;
            11'd7: table_out = 36'heabe4add7;
            11'd8: table_out = 36'heabaab036;
            11'd9: table_out = 36'heab70a978;
            11'd10: table_out = 36'heab36999b;
            11'd11: table_out = 36'heaafc809c;
            11'd12: table_out = 36'heaac25e78;
            11'd13: table_out = 36'heaa88332c;
            11'd14: table_out = 36'heaa4dfeb5;
            11'd15: table_out = 36'heaa13c110;
            11'd16: table_out = 36'hea9d97a3b;
            11'd17: table_out = 36'hea99f2a32;
            11'd18: table_out = 36'hea964d0f3;
            11'd19: table_out = 36'hea92a6e7a;
            11'd20: table_out = 36'hea8f002c6;
            11'd21: table_out = 36'hea8b58dd2;
            11'd22: table_out = 36'hea87b0f9c;
            11'd23: table_out = 36'hea8408821;
            11'd24: table_out = 36'hea805f75e;
            11'd25: table_out = 36'hea7cb5d50;
            11'd26: table_out = 36'hea790b9f4;
            11'd27: table_out = 36'hea7560d48;
            11'd28: table_out = 36'hea71b5748;
            11'd29: table_out = 36'hea6e097f1;
            11'd30: table_out = 36'hea6a5cf40;
            11'd31: table_out = 36'hea66afd32;
            11'd32: table_out = 36'hea63021c5;
            11'd33: table_out = 36'hea5f53cf5;
            11'd34: table_out = 36'hea5ba4ec0;
            11'd35: table_out = 36'hea57f5722;
            11'd36: table_out = 36'hea5445618;
            11'd37: table_out = 36'hea5094b9f;
            11'd38: table_out = 36'hea4ce37b5;
            11'd39: table_out = 36'hea4931a56;
            11'd40: table_out = 36'hea457f380;
            11'd41: table_out = 36'hea41cc32e;
            11'd42: table_out = 36'hea3e1895f;
            11'd43: table_out = 36'hea3a6460f;
            11'd44: table_out = 36'hea36af93b;
            11'd45: table_out = 36'hea32fa2df;
            11'd46: table_out = 36'hea2f442fa;
            11'd47: table_out = 36'hea2b8d988;
            11'd48: table_out = 36'hea27d6686;
            11'd49: table_out = 36'hea241e9f0;
            11'd50: table_out = 36'hea20663c4;
            11'd51: table_out = 36'hea1cad3fe;
            11'd52: table_out = 36'hea18f3a9c;
            11'd53: table_out = 36'hea153979a;
            11'd54: table_out = 36'hea117eaf6;
            11'd55: table_out = 36'hea0dc34ac;
            11'd56: table_out = 36'hea0a074b8;
            11'd57: table_out = 36'hea064ab19;
            11'd58: table_out = 36'hea028d7ca;
            11'd59: table_out = 36'he9fecfac9;
            11'd60: table_out = 36'he9fb11412;
            11'd61: table_out = 36'he9f7523a3;
            11'd62: table_out = 36'he9f392977;
            11'd63: table_out = 36'he9efd258d;
            11'd64: table_out = 36'he9ec117e1;
            11'd65: table_out = 36'he9e85006f;
            11'd66: table_out = 36'he9e48df35;
            11'd67: table_out = 36'he9e0cb42e;
            11'd68: table_out = 36'he9dd07f59;
            11'd69: table_out = 36'he9d9440b2;
            11'd70: table_out = 36'he9d57f836;
            11'd71: table_out = 36'he9d1ba5e1;
            11'd72: table_out = 36'he9cdf49b0;
            11'd73: table_out = 36'he9ca2e3a0;
            11'd74: table_out = 36'he9c6673ae;
            11'd75: table_out = 36'he9c29f9d7;
            11'd76: table_out = 36'he9bed7616;
            11'd77: table_out = 36'he9bb0e86a;
            11'd78: table_out = 36'he9b7450cf;
            11'd79: table_out = 36'he9b37af41;
            11'd80: table_out = 36'he9afb03be;
            11'd81: table_out = 36'he9abe4e41;
            11'd82: table_out = 36'he9a818ec8;
            11'd83: table_out = 36'he9a44c550;
            11'd84: table_out = 36'he9a07f1d5;
            11'd85: table_out = 36'he99cb1453;
            11'd86: table_out = 36'he998e2cc9;
            11'd87: table_out = 36'he99513b31;
            11'd88: table_out = 36'he99143f89;
            11'd89: table_out = 36'he98d739ce;
            11'd90: table_out = 36'he989a29fc;
            11'd91: table_out = 36'he985d1010;
            11'd92: table_out = 36'he981fec06;
            11'd93: table_out = 36'he97e2bddc;
            11'd94: table_out = 36'he97a5858e;
            11'd95: table_out = 36'he97684318;
            11'd96: table_out = 36'he972af677;
            11'd97: table_out = 36'he96ed9fa8;
            11'd98: table_out = 36'he96b03ea7;
            11'd99: table_out = 36'he9672d371;
            11'd100: table_out = 36'he96355e03;
            11'd101: table_out = 36'he95f7de59;
            11'd102: table_out = 36'he95ba5470;
            11'd103: table_out = 36'he957cc044;
            11'd104: table_out = 36'he953f21d1;
            11'd105: table_out = 36'he95017916;
            11'd106: table_out = 36'he94c3c60d;
            11'd107: table_out = 36'he948608b4;
            11'd108: table_out = 36'he94484107;
            11'd109: table_out = 36'he940a6f03;
            11'd110: table_out = 36'he93cc92a4;
            11'd111: table_out = 36'he938eabe7;
            11'd112: table_out = 36'he9350bac8;
            11'd113: table_out = 36'he9312bf44;
            11'd114: table_out = 36'he92d4b958;
            11'd115: table_out = 36'he9296a8ff;
            11'd116: table_out = 36'he92588e36;
            11'd117: table_out = 36'he921a68fa;
            11'd118: table_out = 36'he91dc3947;
            11'd119: table_out = 36'he919dff1a;
            11'd120: table_out = 36'he915fba70;
            11'd121: table_out = 36'he91216b44;
            11'd122: table_out = 36'he90e31193;
            11'd123: table_out = 36'he90a4ad59;
            11'd124: table_out = 36'he90663e94;
            11'd125: table_out = 36'he9027c53f;
            11'd126: table_out = 36'he8fe94157;
            11'd127: table_out = 36'he8faab2d8;
            11'd128: table_out = 36'he8f6c19bf;
            11'd129: table_out = 36'he8f2d7608;
            11'd130: table_out = 36'he8eeec7b0;
            11'd131: table_out = 36'he8eb00eb2;
            11'd132: table_out = 36'he8e714b0c;
            11'd133: table_out = 36'he8e327cb9;
            11'd134: table_out = 36'he8df3a3b6;
            11'd135: table_out = 36'he8db4c000;
            11'd136: table_out = 36'he8d75d192;
            11'd137: table_out = 36'he8d36d86a;
            11'd138: table_out = 36'he8cf7d483;
            11'd139: table_out = 36'he8cb8c5d9;
            11'd140: table_out = 36'he8c79ac6a;
            11'd141: table_out = 36'he8c3a8831;
            11'd142: table_out = 36'he8bfb592b;
            11'd143: table_out = 36'he8bbc1f53;
            11'd144: table_out = 36'he8b7cdaa7;
            11'd145: table_out = 36'he8b3d8b23;
            11'd146: table_out = 36'he8afe30c2;
            11'd147: table_out = 36'he8abecb81;
            11'd148: table_out = 36'he8a7f5b5d;
            11'd149: table_out = 36'he8a3fe052;
            11'd150: table_out = 36'he8a005a5b;
            11'd151: table_out = 36'he89c0c975;
            11'd152: table_out = 36'he89812d9d;
            11'd153: table_out = 36'he894186cf;
            11'd154: table_out = 36'he8901d506;
            11'd155: table_out = 36'he88c2183f;
            11'd156: table_out = 36'he88825077;
            11'd157: table_out = 36'he88427da8;
            11'd158: table_out = 36'he88029fd1;
            11'd159: table_out = 36'he87c2b6ec;
            11'd160: table_out = 36'he8782c2f6;
            11'd161: table_out = 36'he8742c3ec;
            11'd162: table_out = 36'he8702b9c8;
            11'd163: table_out = 36'he86c2a488;
            11'd164: table_out = 36'he86828428;
            11'd165: table_out = 36'he864258a3;
            11'd166: table_out = 36'he860221f6;
            11'd167: table_out = 36'he85c1e01d;
            11'd168: table_out = 36'he85819315;
            11'd169: table_out = 36'he85413ad8;
            11'd170: table_out = 36'he8500d763;
            11'd171: table_out = 36'he84c068b3;
            11'd172: table_out = 36'he847feec4;
            11'd173: table_out = 36'he843f6990;
            11'd174: table_out = 36'he83fed916;
            11'd175: table_out = 36'he83be3d50;
            11'd176: table_out = 36'he837d963a;
            11'd177: table_out = 36'he833ce3d2;
            11'd178: table_out = 36'he82fc2611;
            11'd179: table_out = 36'he82bb5cf6;
            11'd180: table_out = 36'he827a887c;
            11'd181: table_out = 36'he8239a89e;
            11'd182: table_out = 36'he81f8bd59;
            11'd183: table_out = 36'he81b7c6a9;
            11'd184: table_out = 36'he8176c489;
            11'd185: table_out = 36'he8135b6f6;
            11'd186: table_out = 36'he80f49dec;
            11'd187: table_out = 36'he80b37966;
            11'd188: table_out = 36'he80724961;
            11'd189: table_out = 36'he80310dd9;
            11'd190: table_out = 36'he7fefc6c8;
            11'd191: table_out = 36'he7fae742d;
            11'd192: table_out = 36'he7f6d1601;
            11'd193: table_out = 36'he7f2bac42;
            11'd194: table_out = 36'he7eea36ea;
            11'd195: table_out = 36'he7ea8b5f7;
            11'd196: table_out = 36'he7e672963;
            11'd197: table_out = 36'he7e25912c;
            11'd198: table_out = 36'he7de3ed4b;
            11'd199: table_out = 36'he7da23dbe;
            11'd200: table_out = 36'he7d608281;
            11'd201: table_out = 36'he7d1ebb8e;
            11'd202: table_out = 36'he7cdce8e3;
            11'd203: table_out = 36'he7c9b0a7a;
            11'd204: table_out = 36'he7c59204f;
            11'd205: table_out = 36'he7c172a5f;
            11'd206: table_out = 36'he7bd528a5;
            11'd207: table_out = 36'he7b931b1e;
            11'd208: table_out = 36'he7b5101c3;
            11'd209: table_out = 36'he7b0edc93;
            11'd210: table_out = 36'he7accab87;
            11'd211: table_out = 36'he7a8a6e9c;
            11'd212: table_out = 36'he7a4825cf;
            11'd213: table_out = 36'he7a05d119;
            11'd214: table_out = 36'he79c37078;
            11'd215: table_out = 36'he798103e7;
            11'd216: table_out = 36'he793e8b61;
            11'd217: table_out = 36'he78fc06e2;
            11'd218: table_out = 36'he78b97667;
            11'd219: table_out = 36'he7876d9ea;
            11'd220: table_out = 36'he78343167;
            11'd221: table_out = 36'he77f17cda;
            11'd222: table_out = 36'he77aebc3f;
            11'd223: table_out = 36'he776bef91;
            11'd224: table_out = 36'he772916cc;
            11'd225: table_out = 36'he76e631ec;
            11'd226: table_out = 36'he76a340eb;
            11'd227: table_out = 36'he766043c6;
            11'd228: table_out = 36'he761d3a79;
            11'd229: table_out = 36'he75da24fe;
            11'd230: table_out = 36'he75970352;
            11'd231: table_out = 36'he7553d570;
            11'd232: table_out = 36'he75109b54;
            11'd233: table_out = 36'he74cd54f8;
            11'd234: table_out = 36'he748a0259;
            11'd235: table_out = 36'he7446a373;
            11'd236: table_out = 36'he74033840;
            11'd237: table_out = 36'he73bfc0bc;
            11'd238: table_out = 36'he737c3ce3;
            11'd239: table_out = 36'he7338acb0;
            11'd240: table_out = 36'he72f5101f;
            11'd241: table_out = 36'he72b1672b;
            11'd242: table_out = 36'he726db1d0;
            11'd243: table_out = 36'he7229f008;
            11'd244: table_out = 36'he71e621d0;
            11'd245: table_out = 36'he71a24723;
            11'd246: table_out = 36'he715e5ffd;
            11'd247: table_out = 36'he711a6c58;
            11'd248: table_out = 36'he70d66c30;
            11'd249: table_out = 36'he70925f80;
            11'd250: table_out = 36'he704e4645;
            11'd251: table_out = 36'he700a2079;
            11'd252: table_out = 36'he6fc5ee17;
            11'd253: table_out = 36'he6f81af1c;
            11'd254: table_out = 36'he6f3d6382;
            11'd255: table_out = 36'he6ef90b44;
            11'd256: table_out = 36'he6eb4a65e;
            11'd257: table_out = 36'he6e7034cc;
            11'd258: table_out = 36'he6e2bb688;
            11'd259: table_out = 36'he6de72b8e;
            11'd260: table_out = 36'he6da293da;
            11'd261: table_out = 36'he6d5def65;
            11'd262: table_out = 36'he6d193e2d;
            11'd263: table_out = 36'he6cd4802b;
            11'd264: table_out = 36'he6c8fb55b;
            11'd265: table_out = 36'he6c4addb9;
            11'd266: table_out = 36'he6c05f940;
            11'd267: table_out = 36'he6bc107ea;
            11'd268: table_out = 36'he6b7c09b3;
            11'd269: table_out = 36'he6b36fe97;
            11'd270: table_out = 36'he6af1e68f;
            11'd271: table_out = 36'he6aacc199;
            11'd272: table_out = 36'he6a678fae;
            11'd273: table_out = 36'he6a2250c9;
            11'd274: table_out = 36'he69dd04e7;
            11'd275: table_out = 36'he6997ac02;
            11'd276: table_out = 36'he69524615;
            11'd277: table_out = 36'he690cd31b;
            11'd278: table_out = 36'he68c75310;
            11'd279: table_out = 36'he6881c5ee;
            11'd280: table_out = 36'he683c2bb0;
            11'd281: table_out = 36'he67f68452;
            11'd282: table_out = 36'he67b0cfcf;
            11'd283: table_out = 36'he676b0e22;
            11'd284: table_out = 36'he67253f45;
            11'd285: table_out = 36'he66df6333;
            11'd286: table_out = 36'he669979e9;
            11'd287: table_out = 36'he66538360;
            11'd288: table_out = 36'he660d7f94;
            11'd289: table_out = 36'he65c76e7f;
            11'd290: table_out = 36'he6581501d;
            11'd291: table_out = 36'he653b2469;
            11'd292: table_out = 36'he64f4eb5d;
            11'd293: table_out = 36'he64aea4f4;
            11'd294: table_out = 36'he64685129;
            11'd295: table_out = 36'he6421eff8;
            11'd296: table_out = 36'he63db815b;
            11'd297: table_out = 36'he6395054d;
            11'd298: table_out = 36'he634e7bc9;
            11'd299: table_out = 36'he6307e4c9;
            11'd300: table_out = 36'he62c14049;
            11'd301: table_out = 36'he627a8e43;
            11'd302: table_out = 36'he6233ceb2;
            11'd303: table_out = 36'he61ed0192;
            11'd304: table_out = 36'he61a626dc;
            11'd305: table_out = 36'he615f3e8c;
            11'd306: table_out = 36'he6118489c;
            11'd307: table_out = 36'he60d14507;
            11'd308: table_out = 36'he608a33c8;
            11'd309: table_out = 36'he604314d9;
            11'd310: table_out = 36'he5ffbe836;
            11'd311: table_out = 36'he5fb4add9;
            11'd312: table_out = 36'he5f6d65bc;
            11'd313: table_out = 36'he5f260fdb;
            11'd314: table_out = 36'he5edeac30;
            11'd315: table_out = 36'he5e973ab6;
            11'd316: table_out = 36'he5e4fbb67;
            11'd317: table_out = 36'he5e082e3f;
            11'd318: table_out = 36'he5dc09337;
            11'd319: table_out = 36'he5d78ea4a;
            11'd320: table_out = 36'he5d313373;
            11'd321: table_out = 36'he5ce96ead;
            11'd322: table_out = 36'he5ca19bf1;
            11'd323: table_out = 36'he5c59bb3b;
            11'd324: table_out = 36'he5c11cc86;
            11'd325: table_out = 36'he5bc9cfcb;
            11'd326: table_out = 36'he5b81c506;
            11'd327: table_out = 36'he5b39ac30;
            11'd328: table_out = 36'he5af18544;
            11'd329: table_out = 36'he5aa9503e;
            11'd330: table_out = 36'he5a610d16;
            11'd331: table_out = 36'he5a18bbc9;
            11'd332: table_out = 36'he59d05c4f;
            11'd333: table_out = 36'he5987eea4;
            11'd334: table_out = 36'he593f72c2;
            11'd335: table_out = 36'he58f6e8a4;
            11'd336: table_out = 36'he58ae5044;
            11'd337: table_out = 36'he5865a99b;
            11'd338: table_out = 36'he581cf4a6;
            11'd339: table_out = 36'he57d4315d;
            11'd340: table_out = 36'he578b5fbc;
            11'd341: table_out = 36'he57427fbc;
            11'd342: table_out = 36'he56f99159;
            11'd343: table_out = 36'he56b0948c;
            11'd344: table_out = 36'he5667894f;
            11'd345: table_out = 36'he561e6f9d;
            11'd346: table_out = 36'he55d54771;
            11'd347: table_out = 36'he558c10c4;
            11'd348: table_out = 36'he5542cb91;
            11'd349: table_out = 36'he54f977d1;
            11'd350: table_out = 36'he54b01580;
            11'd351: table_out = 36'he5466a497;
            11'd352: table_out = 36'he541d2511;
            11'd353: table_out = 36'he53d396e7;
            11'd354: table_out = 36'he5389fa14;
            11'd355: table_out = 36'he53404e93;
            11'd356: table_out = 36'he52f6945c;
            11'd357: table_out = 36'he52accb6b;
            11'd358: table_out = 36'he5262f3b9;
            11'd359: table_out = 36'he52190d41;
            11'd360: table_out = 36'he51cf17fc;
            11'd361: table_out = 36'he518513e5;
            11'd362: table_out = 36'he513b00f5;
            11'd363: table_out = 36'he50f0df28;
            11'd364: table_out = 36'he50a6ae76;
            11'd365: table_out = 36'he505c6eda;
            11'd366: table_out = 36'he5012204e;
            11'd367: table_out = 36'he4fc7c2cb;
            11'd368: table_out = 36'he4f7d564c;
            11'd369: table_out = 36'he4f32dacb;
            11'd370: table_out = 36'he4ee85042;
            11'd371: table_out = 36'he4e9db6aa;
            11'd372: table_out = 36'he4e530dfe;
            11'd373: table_out = 36'he4e085637;
            11'd374: table_out = 36'he4dbd8f4f;
            11'd375: table_out = 36'he4d72b941;
            11'd376: table_out = 36'he4d27d405;
            11'd377: table_out = 36'he4cdcdf96;
            11'd378: table_out = 36'he4c91dbee;
            11'd379: table_out = 36'he4c46c907;
            11'd380: table_out = 36'he4bfba6d9;
            11'd381: table_out = 36'he4bb07560;
            11'd382: table_out = 36'he4b653494;
            11'd383: table_out = 36'he4b19e470;
            11'd384: table_out = 36'he4ace84ee;
            11'd385: table_out = 36'he4a831606;
            11'd386: table_out = 36'he4a3797b3;
            11'd387: table_out = 36'he49ec09ef;
            11'd388: table_out = 36'he49a06cb2;
            11'd389: table_out = 36'he4954bff8;
            11'd390: table_out = 36'he490903b8;
            11'd391: table_out = 36'he48bd37ee;
            11'd392: table_out = 36'he48715c92;
            11'd393: table_out = 36'he4825719f;
            11'd394: table_out = 36'he47d9770e;
            11'd395: table_out = 36'he478d6cd7;
            11'd396: table_out = 36'he474152f6;
            11'd397: table_out = 36'he46f52964;
            11'd398: table_out = 36'he46a8f019;
            11'd399: table_out = 36'he465ca710;
            11'd400: table_out = 36'he46104e42;
            11'd401: table_out = 36'he45c3e5a8;
            11'd402: table_out = 36'he45776d3c;
            11'd403: table_out = 36'he452ae4f8;
            11'd404: table_out = 36'he44de4cd4;
            11'd405: table_out = 36'he4491a4cb;
            11'd406: table_out = 36'he4444ecd5;
            11'd407: table_out = 36'he43f824ed;
            11'd408: table_out = 36'he43ab4d0b;
            11'd409: table_out = 36'he435e6528;
            11'd410: table_out = 36'he43116d3e;
            11'd411: table_out = 36'he42c46547;
            11'd412: table_out = 36'he42774d3c;
            11'd413: table_out = 36'he422a2515;
            11'd414: table_out = 36'he41dceccd;
            11'd415: table_out = 36'he418fa45c;
            11'd416: table_out = 36'he41424bbb;
            11'd417: table_out = 36'he40f4e2e5;
            11'd418: table_out = 36'he40a769d2;
            11'd419: table_out = 36'he4059e07b;
            11'd420: table_out = 36'he400c46d9;
            11'd421: table_out = 36'he3fbe9ce6;
            11'd422: table_out = 36'he3f70e29b;
            11'd423: table_out = 36'he3f2317f1;
            11'd424: table_out = 36'he3ed53ce0;
            11'd425: table_out = 36'he3e875163;
            11'd426: table_out = 36'he3e395571;
            11'd427: table_out = 36'he3deb4905;
            11'd428: table_out = 36'he3d9d2c17;
            11'd429: table_out = 36'he3d4efea0;
            11'd430: table_out = 36'he3d00c099;
            11'd431: table_out = 36'he3cb271fc;
            11'd432: table_out = 36'he3c6412c0;
            11'd433: table_out = 36'he3c15a2e0;
            11'd434: table_out = 36'he3bc72253;
            11'd435: table_out = 36'he3b789114;
            11'd436: table_out = 36'he3b29ef1a;
            11'd437: table_out = 36'he3adb3c5f;
            11'd438: table_out = 36'he3a8c78db;
            11'd439: table_out = 36'he3a3da487;
            11'd440: table_out = 36'he39eebf5d;
            11'd441: table_out = 36'he399fc955;
            11'd442: table_out = 36'he3950c267;
            11'd443: table_out = 36'he3901aa8d;
            11'd444: table_out = 36'he38b281bf;
            11'd445: table_out = 36'he386347f6;
            11'd446: table_out = 36'he3813fd2a;
            11'd447: table_out = 36'he37c4a155;
            11'd448: table_out = 36'he37753470;
            11'd449: table_out = 36'he3725b671;
            11'd450: table_out = 36'he36d62753;
            11'd451: table_out = 36'he3686870e;
            11'd452: table_out = 36'he3636d59b;
            11'd453: table_out = 36'he35e712f1;
            11'd454: table_out = 36'he35973f0b;
            11'd455: table_out = 36'he354759df;
            11'd456: table_out = 36'he34f76367;
            11'd457: table_out = 36'he34a75b9c;
            11'd458: table_out = 36'he34574275;
            11'd459: table_out = 36'he340717eb;
            11'd460: table_out = 36'he33b6dbf7;
            11'd461: table_out = 36'he33668e91;
            11'd462: table_out = 36'he33162fb2;
            11'd463: table_out = 36'he32c5bf51;
            11'd464: table_out = 36'he32753d68;
            11'd465: table_out = 36'he3224a9ee;
            11'd466: table_out = 36'he31d404dc;
            11'd467: table_out = 36'he31834e2a;
            11'd468: table_out = 36'he313285d1;
            11'd469: table_out = 36'he30e1abc9;
            11'd470: table_out = 36'he3090c009;
            11'd471: table_out = 36'he303fc28b;
            11'd472: table_out = 36'he2feeb346;
            11'd473: table_out = 36'he2f9d9233;
            11'd474: table_out = 36'he2f4c5f4a;
            11'd475: table_out = 36'he2efb1a82;
            11'd476: table_out = 36'he2ea9c3d5;
            11'd477: table_out = 36'he2e585b3a;
            11'd478: table_out = 36'he2e06e0aa;
            11'd479: table_out = 36'he2db5541b;
            11'd480: table_out = 36'he2d63b587;
            11'd481: table_out = 36'he2d1204e6;
            11'd482: table_out = 36'he2cc0422f;
            11'd483: table_out = 36'he2c6e6d5b;
            11'd484: table_out = 36'he2c1c8660;
            11'd485: table_out = 36'he2bca8d39;
            11'd486: table_out = 36'he2b7881db;
            11'd487: table_out = 36'he2b266440;
            11'd488: table_out = 36'he2ad4345f;
            11'd489: table_out = 36'he2a81f22f;
            11'd490: table_out = 36'he2a2f9daa;
            11'd491: table_out = 36'he29dd36c6;
            11'd492: table_out = 36'he298abd7b;
            11'd493: table_out = 36'he293831c2;
            11'd494: table_out = 36'he28e59391;
            11'd495: table_out = 36'he2892e2e1;
            11'd496: table_out = 36'he28401fa9;
            11'd497: table_out = 36'he27ed49e2;
            11'd498: table_out = 36'he279a6182;
            11'd499: table_out = 36'he27476681;
            11'd500: table_out = 36'he26f458d8;
            11'd501: table_out = 36'he26a1387d;
            11'd502: table_out = 36'he264e0568;
            11'd503: table_out = 36'he25fabf91;
            11'd504: table_out = 36'he25a766ef;
            11'd505: table_out = 36'he2553fb79;
            11'd506: table_out = 36'he25007d28;
            11'd507: table_out = 36'he24acebf3;
            11'd508: table_out = 36'he245947d1;
            11'd509: table_out = 36'he240590b9;
            11'd510: table_out = 36'he23b1c6a4;
            11'd511: table_out = 36'he235de987;
            11'd512: table_out = 36'he2309f95c;
            11'd513: table_out = 36'he22b5f618;
            11'd514: table_out = 36'he2261dfb4;
            11'd515: table_out = 36'he220db626;
            11'd516: table_out = 36'he21b97966;
            11'd517: table_out = 36'he2165296c;
            11'd518: table_out = 36'he2110c62d;
            11'd519: table_out = 36'he20bc4fa2;
            11'd520: table_out = 36'he2067c5c2;
            11'd521: table_out = 36'he20132883;
            11'd522: table_out = 36'he1fbe77de;
            11'd523: table_out = 36'he1f69b3c8;
            11'd524: table_out = 36'he1f14dc3a;
            11'd525: table_out = 36'he1ebff129;
            11'd526: table_out = 36'he1e6af28e;
            11'd527: table_out = 36'he1e15e05f;
            11'd528: table_out = 36'he1dc0ba93;
            11'd529: table_out = 36'he1d6b8121;
            11'd530: table_out = 36'he1d163400;
            11'd531: table_out = 36'he1cc0d328;
            11'd532: table_out = 36'he1c6b5e8d;
            11'd533: table_out = 36'he1c15d629;
            11'd534: table_out = 36'he1bc039f1;
            11'd535: table_out = 36'he1b6a89dc;
            11'd536: table_out = 36'he1b14c5e1;
            11'd537: table_out = 36'he1abeedf7;
            11'd538: table_out = 36'he1a690214;
            11'd539: table_out = 36'he1a130230;
            11'd540: table_out = 36'he19bcee40;
            11'd541: table_out = 36'he1966c63c;
            11'd542: table_out = 36'he19108a1a;
            11'd543: table_out = 36'he18ba39d1;
            11'd544: table_out = 36'he1863d557;
            11'd545: table_out = 36'he180d5ca3;
            11'd546: table_out = 36'he17b6cfab;
            11'd547: table_out = 36'he17602e66;
            11'd548: table_out = 36'he170978cb;
            11'd549: table_out = 36'he16b2aecf;
            11'd550: table_out = 36'he165bd06a;
            11'd551: table_out = 36'he1604dd91;
            11'd552: table_out = 36'he15add63b;
            11'd553: table_out = 36'he1556ba5e;
            11'd554: table_out = 36'he14ff89f1;
            11'd555: table_out = 36'he14a844ea;
            11'd556: table_out = 36'he1450eb3f;
            11'd557: table_out = 36'he13f97ce6;
            11'd558: table_out = 36'he13a1f9d6;
            11'd559: table_out = 36'he134a6204;
            11'd560: table_out = 36'he12f2b567;
            11'd561: table_out = 36'he129af3f6;
            11'd562: table_out = 36'he12431da5;
            11'd563: table_out = 36'he11eb326c;
            11'd564: table_out = 36'he1193323f;
            11'd565: table_out = 36'he113b1d16;
            11'd566: table_out = 36'he10e2f2e6;
            11'd567: table_out = 36'he108ab3a6;
            11'd568: table_out = 36'he10325f4a;
            11'd569: table_out = 36'he0fd9f5c9;
            11'd570: table_out = 36'he0f817719;
            11'd571: table_out = 36'he0f28e330;
            11'd572: table_out = 36'he0ed03a03;
            11'd573: table_out = 36'he0e777b88;
            11'd574: table_out = 36'he0e1ea7b5;
            11'd575: table_out = 36'he0dc5be80;
            11'd576: table_out = 36'he0d6cbfdf;
            11'd577: table_out = 36'he0d13abc6;
            11'd578: table_out = 36'he0cba822c;
            11'd579: table_out = 36'he0c614307;
            11'd580: table_out = 36'he0c07ee4b;
            11'd581: table_out = 36'he0bae83ef;
            11'd582: table_out = 36'he0b5503e8;
            11'd583: table_out = 36'he0afb6e2b;
            11'd584: table_out = 36'he0aa1c2ae;
            11'd585: table_out = 36'he0a480166;
            11'd586: table_out = 36'he09ee2a49;
            11'd587: table_out = 36'he09943d4d;
            11'd588: table_out = 36'he093a3a65;
            11'd589: table_out = 36'he08e02189;
            11'd590: table_out = 36'he0885f2ac;
            11'd591: table_out = 36'he082badc5;
            11'd592: table_out = 36'he07d152c8;
            11'd593: table_out = 36'he0776e1ab;
            11'd594: table_out = 36'he071c5a63;
            11'd595: table_out = 36'he06c1bce4;
            11'd596: table_out = 36'he06670925;
            11'd597: table_out = 36'he060c3f19;
            11'd598: table_out = 36'he05b15eb7;
            11'd599: table_out = 36'he055667f3;
            11'd600: table_out = 36'he04fb5ac2;
            11'd601: table_out = 36'he04a03719;
            11'd602: table_out = 36'he0444fced;
            11'd603: table_out = 36'he03e9ac33;
            11'd604: table_out = 36'he038e44df;
            11'd605: table_out = 36'he0332c6e7;
            11'd606: table_out = 36'he02d7323f;
            11'd607: table_out = 36'he027b86db;
            11'd608: table_out = 36'he021fc4b2;
            11'd609: table_out = 36'he01c3ebb7;
            11'd610: table_out = 36'he0167fbde;
            11'd611: table_out = 36'he010bf51d;
            11'd612: table_out = 36'he00afd769;
            11'd613: table_out = 36'he0053a2b5;
            11'd614: table_out = 36'hdfff756f6;
            11'd615: table_out = 36'hdff9af421;
            11'd616: table_out = 36'hdff3e7a2a;
            11'd617: table_out = 36'hdfee1e905;
            11'd618: table_out = 36'hdfe8540a7;
            11'd619: table_out = 36'hdfe288104;
            11'd620: table_out = 36'hdfdcbaa11;
            11'd621: table_out = 36'hdfd6ebbc2;
            11'd622: table_out = 36'hdfd11b60b;
            11'd623: table_out = 36'hdfcb498df;
            11'd624: table_out = 36'hdfc576434;
            11'd625: table_out = 36'hdfbfa17fe;
            11'd626: table_out = 36'hdfb9cb430;
            11'd627: table_out = 36'hdfb3f38bf;
            11'd628: table_out = 36'hdfae1a59e;
            11'd629: table_out = 36'hdfa83fac2;
            11'd630: table_out = 36'hdfa26381f;
            11'd631: table_out = 36'hdf9c85da8;
            11'd632: table_out = 36'hdf96a6b52;
            11'd633: table_out = 36'hdf90c6110;
            11'd634: table_out = 36'hdf8ae3ed5;
            11'd635: table_out = 36'hdf8500497;
            11'd636: table_out = 36'hdf7f1b248;
            11'd637: table_out = 36'hdf79347dc;
            11'd638: table_out = 36'hdf734c547;
            11'd639: table_out = 36'hdf6d62a7d;
            11'd640: table_out = 36'hdf6777771;
            11'd641: table_out = 36'hdf618ac16;
            11'd642: table_out = 36'hdf5b9c861;
            11'd643: table_out = 36'hdf55acc44;
            11'd644: table_out = 36'hdf4fbb7b3;
            11'd645: table_out = 36'hdf49c8aa2;
            11'd646: table_out = 36'hdf43d4504;
            11'd647: table_out = 36'hdf3dde6cb;
            11'd648: table_out = 36'hdf37e6fec;
            11'd649: table_out = 36'hdf31ee05a;
            11'd650: table_out = 36'hdf2bf3808;
            11'd651: table_out = 36'hdf25f76e8;
            11'd652: table_out = 36'hdf1ff9cef;
            11'd653: table_out = 36'hdf19faa0f;
            11'd654: table_out = 36'hdf13f9e3b;
            11'd655: table_out = 36'hdf0df7967;
            11'd656: table_out = 36'hdf07f3b85;
            11'd657: table_out = 36'hdf01ee488;
            11'd658: table_out = 36'hdefbe7463;
            11'd659: table_out = 36'hdef5deb09;
            11'd660: table_out = 36'hdeefd486d;
            11'd661: table_out = 36'hdee9c8c81;
            11'd662: table_out = 36'hdee3bb739;
            11'd663: table_out = 36'hdeddac887;
            11'd664: table_out = 36'hded79c05d;
            11'd665: table_out = 36'hded189eae;
            11'd666: table_out = 36'hdecb7636d;
            11'd667: table_out = 36'hdec560e8d;
            11'd668: table_out = 36'hdebf49fff;
            11'd669: table_out = 36'hdeb9317b6;
            11'd670: table_out = 36'hdeb3175a5;
            11'd671: table_out = 36'hdeacfb9be;
            11'd672: table_out = 36'hdea6de3f3;
            11'd673: table_out = 36'hdea0bf436;
            11'd674: table_out = 36'hde9a9ea7b;
            11'd675: table_out = 36'hde947c6b2;
            11'd676: table_out = 36'hde8e588ce;
            11'd677: table_out = 36'hde88330c2;
            11'd678: table_out = 36'hde820be7e;
            11'd679: table_out = 36'hde7be31f6;
            11'd680: table_out = 36'hde75b8b1c;
            11'd681: table_out = 36'hde6f8c9e0;
            11'd682: table_out = 36'hde695ee35;
            11'd683: table_out = 36'hde632f80d;
            11'd684: table_out = 36'hde5cfe75a;
            11'd685: table_out = 36'hde56cbc0d;
            11'd686: table_out = 36'hde5097618;
            11'd687: table_out = 36'hde4a6156d;
            11'd688: table_out = 36'hde44299fe;
            11'd689: table_out = 36'hde3df03bb;
            11'd690: table_out = 36'hde37b5296;
            11'd691: table_out = 36'hde3178682;
            11'd692: table_out = 36'hde2b39f6f;
            11'd693: table_out = 36'hde24f9d4e;
            11'd694: table_out = 36'hde1eb8012;
            11'd695: table_out = 36'hde18747aa;
            11'd696: table_out = 36'hde122f40a;
            11'd697: table_out = 36'hde0be8521;
            11'd698: table_out = 36'hde059fae1;
            11'd699: table_out = 36'hddff5553b;
            11'd700: table_out = 36'hddf909420;
            11'd701: table_out = 36'hddf2bb782;
            11'd702: table_out = 36'hddec6bf50;
            11'd703: table_out = 36'hdde61ab7c;
            11'd704: table_out = 36'hdddfc7bf7;
            11'd705: table_out = 36'hddd9730b1;
            11'd706: table_out = 36'hddd31c99c;
            11'd707: table_out = 36'hddccc46a8;
            11'd708: table_out = 36'hddc66a7c6;
            11'd709: table_out = 36'hddc00ece5;
            11'd710: table_out = 36'hddb9b15f8;
            11'd711: table_out = 36'hddb3522ef;
            11'd712: table_out = 36'hddacf13b9;
            11'd713: table_out = 36'hdda68e847;
            11'd714: table_out = 36'hdda02a08a;
            11'd715: table_out = 36'hdd99c3c72;
            11'd716: table_out = 36'hdd935bbf0;
            11'd717: table_out = 36'hdd8cf1ef2;
            11'd718: table_out = 36'hdd868656b;
            11'd719: table_out = 36'hdd8018f49;
            11'd720: table_out = 36'hdd79a9c7c;
            11'd721: table_out = 36'hdd7338cf6;
            11'd722: table_out = 36'hdd6cc60a5;
            11'd723: table_out = 36'hdd665177a;
            11'd724: table_out = 36'hdd5fdb164;
            11'd725: table_out = 36'hdd5962e53;
            11'd726: table_out = 36'hdd52e8e38;
            11'd727: table_out = 36'hdd4c6d101;
            11'd728: table_out = 36'hdd45ef69e;
            11'd729: table_out = 36'hdd3f6ff00;
            11'd730: table_out = 36'hdd38eea14;
            11'd731: table_out = 36'hdd326b7cc;
            11'd732: table_out = 36'hdd2be6816;
            11'd733: table_out = 36'hdd255fae1;
            11'd734: table_out = 36'hdd1ed701e;
            11'd735: table_out = 36'hdd184c7ba;
            11'd736: table_out = 36'hdd11c01a6;
            11'd737: table_out = 36'hdd0b31dd0;
            11'd738: table_out = 36'hdd04a1c28;
            11'd739: table_out = 36'hdcfe0fc9d;
            11'd740: table_out = 36'hdcf77bf1d;
            11'd741: table_out = 36'hdcf0e6398;
            11'd742: table_out = 36'hdcea4e9fc;
            11'd743: table_out = 36'hdce3b5238;
            11'd744: table_out = 36'hdcdd19c3b;
            11'd745: table_out = 36'hdcd67c7f4;
            11'd746: table_out = 36'hdccfdd550;
            11'd747: table_out = 36'hdcc93c440;
            11'd748: table_out = 36'hdcc2994b1;
            11'd749: table_out = 36'hdcbbf4691;
            11'd750: table_out = 36'hdcb54d9d0;
            11'd751: table_out = 36'hdcaea4e5a;
            11'd752: table_out = 36'hdca7fa420;
            11'd753: table_out = 36'hdca14db0e;
            11'd754: table_out = 36'hdc9a9f314;
            11'd755: table_out = 36'hdc93eec1e;
            11'd756: table_out = 36'hdc8d3c61c;
            11'd757: table_out = 36'hdc86880fb;
            11'd758: table_out = 36'hdc7fd1ca9;
            11'd759: table_out = 36'hdc7919913;
            11'd760: table_out = 36'hdc725f628;
            11'd761: table_out = 36'hdc6ba33d6;
            11'd762: table_out = 36'hdc64e5209;
            11'd763: table_out = 36'hdc5e250b0;
            11'd764: table_out = 36'hdc5762fb8;
            11'd765: table_out = 36'hdc509ef0f;
            11'd766: table_out = 36'hdc49d8ea2;
            11'd767: table_out = 36'hdc4310e5e;
            11'd768: table_out = 36'hdc3c46e30;
            11'd769: table_out = 36'hdc357ae07;
            11'd770: table_out = 36'hdc2eacdce;
            11'd771: table_out = 36'hdc27dcd73;
            11'd772: table_out = 36'hdc210ace3;
            11'd773: table_out = 36'hdc1a36c0b;
            11'd774: table_out = 36'hdc1360ad8;
            11'd775: table_out = 36'hdc0c88937;
            11'd776: table_out = 36'hdc05ae714;
            11'd777: table_out = 36'hdbfed245c;
            11'd778: table_out = 36'hdbf7f40fc;
            11'd779: table_out = 36'hdbf113ce0;
            11'd780: table_out = 36'hdbea317f4;
            11'd781: table_out = 36'hdbe34d226;
            11'd782: table_out = 36'hdbdc66b61;
            11'd783: table_out = 36'hdbd57e392;
            11'd784: table_out = 36'hdbce93aa5;
            11'd785: table_out = 36'hdbc7a7086;
            11'd786: table_out = 36'hdbc0b8521;
            11'd787: table_out = 36'hdbb9c7862;
            11'd788: table_out = 36'hdbb2d4a35;
            11'd789: table_out = 36'hdbabdfa86;
            11'd790: table_out = 36'hdba4e8940;
            11'd791: table_out = 36'hdb9def650;
            11'd792: table_out = 36'hdb96f41a1;
            11'd793: table_out = 36'hdb8ff6b1f;
            11'd794: table_out = 36'hdb88f72b4;
            11'd795: table_out = 36'hdb81f584d;
            11'd796: table_out = 36'hdb7af1bd5;
            11'd797: table_out = 36'hdb73ebd37;
            11'd798: table_out = 36'hdb6ce3c5e;
            11'd799: table_out = 36'hdb65d9936;
            11'd800: table_out = 36'hdb5ecd3a8;
            11'd801: table_out = 36'hdb57beba2;
            11'd802: table_out = 36'hdb50ae10c;
            11'd803: table_out = 36'hdb499b3d3;
            11'd804: table_out = 36'hdb42863e1;
            11'd805: table_out = 36'hdb3b6f120;
            11'd806: table_out = 36'hdb3455b7b;
            11'd807: table_out = 36'hdb2d3a2dd;
            11'd808: table_out = 36'hdb261c730;
            11'd809: table_out = 36'hdb1efc85f;
            11'd810: table_out = 36'hdb17da653;
            11'd811: table_out = 36'hdb10b60f7;
            11'd812: table_out = 36'hdb098f835;
            11'd813: table_out = 36'hdb0266bf7;
            11'd814: table_out = 36'hdafb3bc27;
            11'd815: table_out = 36'hdaf40e8af;
            11'd816: table_out = 36'hdaecdf179;
            11'd817: table_out = 36'hdae5ad66f;
            11'd818: table_out = 36'hdade79779;
            11'd819: table_out = 36'hdad743482;
            11'd820: table_out = 36'hdad00ad73;
            11'd821: table_out = 36'hdac8d0236;
            11'd822: table_out = 36'hdac1932b3;
            11'd823: table_out = 36'hdaba53ed5;
            11'd824: table_out = 36'hdab312683;
            11'd825: table_out = 36'hdaabce9a8;
            11'd826: table_out = 36'hdaa48882d;
            11'd827: table_out = 36'hda9d401f9;
            11'd828: table_out = 36'hda95f56f6;
            11'd829: table_out = 36'hda8ea870d;
            11'd830: table_out = 36'hda8759226;
            11'd831: table_out = 36'hda800782a;
            11'd832: table_out = 36'hda78b3901;
            11'd833: table_out = 36'hda715d493;
            11'd834: table_out = 36'hda6a04aca;
            11'd835: table_out = 36'hda62a9b8d;
            11'd836: table_out = 36'hda5b4c6c3;
            11'd837: table_out = 36'hda53ecc57;
            11'd838: table_out = 36'hda4c8ac2e;
            11'd839: table_out = 36'hda4526631;
            11'd840: table_out = 36'hda3dbfa48;
            11'd841: table_out = 36'hda365685a;
            11'd842: table_out = 36'hda2eeb04f;
            11'd843: table_out = 36'hda277d20e;
            11'd844: table_out = 36'hda200cd80;
            11'd845: table_out = 36'hda189a28a;
            11'd846: table_out = 36'hda1125114;
            11'd847: table_out = 36'hda09ad906;
            11'd848: table_out = 36'hda0233a46;
            11'd849: table_out = 36'hd9fab74bc;
            11'd850: table_out = 36'hd9f33884d;
            11'd851: table_out = 36'hd9ebb74e1;
            11'd852: table_out = 36'hd9e433a5e;
            11'd853: table_out = 36'hd9dcad8ab;
            11'd854: table_out = 36'hd9d524faf;
            11'd855: table_out = 36'hd9cd99f4f;
            11'd856: table_out = 36'hd9c60c772;
            11'd857: table_out = 36'hd9be7c7fe;
            11'd858: table_out = 36'hd9b6ea0d9;
            11'd859: table_out = 36'hd9af551e9;
            11'd860: table_out = 36'hd9a7bdb13;
            11'd861: table_out = 36'hd9a023c3e;
            11'd862: table_out = 36'hd9988754f;
            11'd863: table_out = 36'hd990e862c;
            11'd864: table_out = 36'hd98946eba;
            11'd865: table_out = 36'hd981a2ede;
            11'd866: table_out = 36'hd979fc67d;
            11'd867: table_out = 36'hd9725357e;
            11'd868: table_out = 36'hd96aa7bc4;
            11'd869: table_out = 36'hd962f9934;
            11'd870: table_out = 36'hd95b48db4;
            11'd871: table_out = 36'hd95395928;
            11'd872: table_out = 36'hd94bdfb74;
            11'd873: table_out = 36'hd9442747e;
            11'd874: table_out = 36'hd93c6c429;
            11'd875: table_out = 36'hd934aea5a;
            11'd876: table_out = 36'hd92cee6f4;
            11'd877: table_out = 36'hd9252b9dd;
            11'd878: table_out = 36'hd91d662f7;
            11'd879: table_out = 36'hd9159e227;
            11'd880: table_out = 36'hd90dd3750;
            11'd881: table_out = 36'hd90606256;
            11'd882: table_out = 36'hd8fe3631d;
            11'd883: table_out = 36'hd8f663987;
            11'd884: table_out = 36'hd8ee8e578;
            11'd885: table_out = 36'hd8e6b66d4;
            11'd886: table_out = 36'hd8dedbd7d;
            11'd887: table_out = 36'hd8d6fe955;
            11'd888: table_out = 36'hd8cf1ea41;
            11'd889: table_out = 36'hd8c73c022;
            11'd890: table_out = 36'hd8bf56adb;
            11'd891: table_out = 36'hd8b76ea4f;
            11'd892: table_out = 36'hd8af83e5f;
            11'd893: table_out = 36'hd8a7966ef;
            11'd894: table_out = 36'hd89fa63e0;
            11'd895: table_out = 36'hd897b3514;
            11'd896: table_out = 36'hd88fbda6c;
            11'd897: table_out = 36'hd887c53cc;
            11'd898: table_out = 36'hd87fca113;
            11'd899: table_out = 36'hd877cc225;
            11'd900: table_out = 36'hd86fcb6e1;
            11'd901: table_out = 36'hd867c7f2a;
            11'd902: table_out = 36'hd85fc1adf;
            11'd903: table_out = 36'hd857b89e4;
            11'd904: table_out = 36'hd84facc17;
            11'd905: table_out = 36'hd8479e15a;
            11'd906: table_out = 36'hd83f8c98e;
            11'd907: table_out = 36'hd83778493;
            11'd908: table_out = 36'hd82f61248;
            11'd909: table_out = 36'hd82747290;
            11'd910: table_out = 36'hd81f2a549;
            11'd911: table_out = 36'hd8170aa53;
            11'd912: table_out = 36'hd80ee818e;
            11'd913: table_out = 36'hd806c2adb;
            11'd914: table_out = 36'hd7fe9a617;
            11'd915: table_out = 36'hd7f66f324;
            11'd916: table_out = 36'hd7ee411e0;
            11'd917: table_out = 36'hd7e61022a;
            11'd918: table_out = 36'hd7dddc3e1;
            11'd919: table_out = 36'hd7d5a56e4;
            11'd920: table_out = 36'hd7cd6bb12;
            11'd921: table_out = 36'hd7c52f04a;
            11'd922: table_out = 36'hd7bcef669;
            11'd923: table_out = 36'hd7b4acd4e;
            11'd924: table_out = 36'hd7ac674d8;
            11'd925: table_out = 36'hd7a41ece4;
            11'd926: table_out = 36'hd79bd3550;
            11'd927: table_out = 36'hd79384df9;
            11'd928: table_out = 36'hd78b336bf;
            11'd929: table_out = 36'hd782def7d;
            11'd930: table_out = 36'hd77a87811;
            11'd931: table_out = 36'hd7722d059;
            11'd932: table_out = 36'hd769cf831;
            11'd933: table_out = 36'hd7616ef76;
            11'd934: table_out = 36'hd7590b605;
            11'd935: table_out = 36'hd750a4bba;
            11'd936: table_out = 36'hd7483b072;
            11'd937: table_out = 36'hd73fce409;
            11'd938: table_out = 36'hd7375e65b;
            11'd939: table_out = 36'hd72eeb744;
            11'd940: table_out = 36'hd726756a0;
            11'd941: table_out = 36'hd71dfc44a;
            11'd942: table_out = 36'hd7158001f;
            11'd943: table_out = 36'hd70d009f8;
            11'd944: table_out = 36'hd7047e1b2;
            11'd945: table_out = 36'hd6fbf8727;
            11'd946: table_out = 36'hd6f36fa32;
            11'd947: table_out = 36'hd6eae3aaf;
            11'd948: table_out = 36'hd6e254876;
            11'd949: table_out = 36'hd6d9c2363;
            11'd950: table_out = 36'hd6d12cb50;
            11'd951: table_out = 36'hd6c894017;
            11'd952: table_out = 36'hd6bff8192;
            11'd953: table_out = 36'hd6b758f9a;
            11'd954: table_out = 36'hd6aeb6a09;
            11'd955: table_out = 36'hd6a6110b8;
            11'd956: table_out = 36'hd69d68380;
            11'd957: table_out = 36'hd694bc23b;
            11'd958: table_out = 36'hd68c0ccc2;
            11'd959: table_out = 36'hd6835a2ec;
            11'd960: table_out = 36'hd67aa4492;
            11'd961: table_out = 36'hd671eb18e;
            11'd962: table_out = 36'hd6692e9b6;
            11'd963: table_out = 36'hd6606ece3;
            11'd964: table_out = 36'hd657abaec;
            11'd965: table_out = 36'hd64ee53aa;
            11'd966: table_out = 36'hd6461b6f3;
            11'd967: table_out = 36'hd63d4e4a0;
            11'd968: table_out = 36'hd6347dc86;
            11'd969: table_out = 36'hd62ba9e7c;
            11'd970: table_out = 36'hd622d2a5b;
            11'd971: table_out = 36'hd619f7ff7;
            11'd972: table_out = 36'hd61119f27;
            11'd973: table_out = 36'hd608387c2;
            11'd974: table_out = 36'hd5ff5399d;
            11'd975: table_out = 36'hd5f66b48e;
            11'd976: table_out = 36'hd5ed7f86b;
            11'd977: table_out = 36'hd5e490509;
            11'd978: table_out = 36'hd5db9da3d;
            11'd979: table_out = 36'hd5d2a77dc;
            11'd980: table_out = 36'hd5c9addbb;
            11'd981: table_out = 36'hd5c0b0bae;
            11'd982: table_out = 36'hd5b7b018a;
            11'd983: table_out = 36'hd5aeabf24;
            11'd984: table_out = 36'hd5a5a444e;
            11'd985: table_out = 36'hd59c990dd;
            11'd986: table_out = 36'hd5938a4a5;
            11'd987: table_out = 36'hd58a77f78;
            11'd988: table_out = 36'hd5816212a;
            11'd989: table_out = 36'hd5784898e;
            11'd990: table_out = 36'hd56f2b877;
            11'd991: table_out = 36'hd5660adb7;
            11'd992: table_out = 36'hd55ce6920;
            11'd993: table_out = 36'hd553bea85;
            11'd994: table_out = 36'hd54a931b8;
            11'd995: table_out = 36'hd54163e89;
            11'd996: table_out = 36'hd538310cc;
            11'd997: table_out = 36'hd52efa850;
            11'd998: table_out = 36'hd525c04e7;
            11'd999: table_out = 36'hd51c82663;
            11'd1000: table_out = 36'hd51340c92;
            11'd1001: table_out = 36'hd509fb746;
            11'd1002: table_out = 36'hd500b264f;
            11'd1003: table_out = 36'hd4f76597d;
            11'd1004: table_out = 36'hd4ee150a0;
            11'd1005: table_out = 36'hd4e4c0b86;
            11'd1006: table_out = 36'hd4db68a00;
            11'd1007: table_out = 36'hd4d20cbdb;
            11'd1008: table_out = 36'hd4c8ad0e8;
            11'd1009: table_out = 36'hd4bf498f5;
            11'd1010: table_out = 36'hd4b5e23cf;
            11'd1011: table_out = 36'hd4ac77145;
            11'd1012: table_out = 36'hd4a308124;
            11'd1013: table_out = 36'hd4999533b;
            11'd1014: table_out = 36'hd4901e757;
            11'd1015: table_out = 36'hd486a3d44;
            11'd1016: table_out = 36'hd47d254d0;
            11'd1017: table_out = 36'hd473a2dc7;
            11'd1018: table_out = 36'hd46a1c7f5;
            11'd1019: table_out = 36'hd46092328;
            11'd1020: table_out = 36'hd45703f29;
            11'd1021: table_out = 36'hd44d71bc6;
            11'd1022: table_out = 36'hd443db8c9;
            11'd1023: table_out = 36'hd43a415fd;
            11'd1024: table_out = 36'hd430a332e;
            11'd1025: table_out = 36'hd42701026;
            11'd1026: table_out = 36'hd41d5acaf;
            11'd1027: table_out = 36'hd413b0893;
            11'd1028: table_out = 36'hd40a0239c;
            11'd1029: table_out = 36'hd4004fd94;
            11'd1030: table_out = 36'hd3f699643;
            11'd1031: table_out = 36'hd3ecded74;
            11'd1032: table_out = 36'hd3e3202ed;
            11'd1033: table_out = 36'hd3d95d679;
            11'd1034: table_out = 36'hd3cf967de;
            11'd1035: table_out = 36'hd3c5cb6e6;
            11'd1036: table_out = 36'hd3bbfc357;
            11'd1037: table_out = 36'hd3b228cf8;
            11'd1038: table_out = 36'hd3a851392;
            11'd1039: table_out = 36'hd39e756ea;
            11'd1040: table_out = 36'hd394956c7;
            11'd1041: table_out = 36'hd38ab12ef;
            11'd1042: table_out = 36'hd380c8b29;
            11'd1043: table_out = 36'hd376dbf39;
            11'd1044: table_out = 36'hd36ceaee5;
            11'd1045: table_out = 36'hd362f59f1;
            11'd1046: table_out = 36'hd358fc024;
            11'd1047: table_out = 36'hd34efe140;
            11'd1048: table_out = 36'hd344fbd0b;
            11'd1049: table_out = 36'hd33af5347;
            11'd1050: table_out = 36'hd330ea3b9;
            11'd1051: table_out = 36'hd326dae24;
            11'd1052: table_out = 36'hd31cc7249;
            11'd1053: table_out = 36'hd312aefed;
            11'd1054: table_out = 36'hd308926d1;
            11'd1055: table_out = 36'hd2fe716b6;
            11'd1056: table_out = 36'hd2f44bf60;
            11'd1057: table_out = 36'hd2ea2208e;
            11'd1058: table_out = 36'hd2dff3a03;
            11'd1059: table_out = 36'hd2d5c0b7d;
            11'd1060: table_out = 36'hd2cb894bf;
            11'd1061: table_out = 36'hd2c14d587;
            11'd1062: table_out = 36'hd2b70cd96;
            11'd1063: table_out = 36'hd2acc7caa;
            11'd1064: table_out = 36'hd2a27e283;
            11'd1065: table_out = 36'hd2982fedf;
            11'd1066: table_out = 36'hd28ddd17c;
            11'd1067: table_out = 36'hd28385a19;
            11'd1068: table_out = 36'hd27929873;
            11'd1069: table_out = 36'hd26ec8c47;
            11'd1070: table_out = 36'hd26463552;
            11'd1071: table_out = 36'hd259f9350;
            11'd1072: table_out = 36'hd24f8a5ff;
            11'd1073: table_out = 36'hd24516d19;
            11'd1074: table_out = 36'hd23a9e85a;
            11'd1075: table_out = 36'hd2302177d;
            11'd1076: table_out = 36'hd2259fa3c;
            11'd1077: table_out = 36'hd21b19053;
            11'd1078: table_out = 36'hd2108d97b;
            11'd1079: table_out = 36'hd205fd56d;
            11'd1080: table_out = 36'hd1fb683e4;
            11'd1081: table_out = 36'hd1f0ce497;
            11'd1082: table_out = 36'hd1e62f73f;
            11'd1083: table_out = 36'hd1db8bb94;
            11'd1084: table_out = 36'hd1d0e314e;
            11'd1085: table_out = 36'hd1c635824;
            11'd1086: table_out = 36'hd1bb82fce;
            11'd1087: table_out = 36'hd1b0cb800;
            11'd1088: table_out = 36'hd1a60f072;
            11'd1089: table_out = 36'hd19b4d8da;
            11'd1090: table_out = 36'hd190870ec;
            11'd1091: table_out = 36'hd185bb85d;
            11'd1092: table_out = 36'hd17aeaee2;
            11'd1093: table_out = 36'hd1701542f;
            11'd1094: table_out = 36'hd1653a7f8;
            11'd1095: table_out = 36'hd15a5a9ef;
            11'd1096: table_out = 36'hd14f759c8;
            11'd1097: table_out = 36'hd1448b734;
            11'd1098: table_out = 36'hd1399c1e6;
            11'd1099: table_out = 36'hd12ea798f;
            11'd1100: table_out = 36'hd123adde1;
            11'd1101: table_out = 36'hd118aee8b;
            11'd1102: table_out = 36'hd10daab3e;
            11'd1103: table_out = 36'hd102a13aa;
            11'd1104: table_out = 36'hd0f79277d;
            11'd1105: table_out = 36'hd0ec7e668;
            11'd1106: table_out = 36'hd0e165017;
            11'd1107: table_out = 36'hd0d64643a;
            11'd1108: table_out = 36'hd0cb2227c;
            11'd1109: table_out = 36'hd0bff8a8c;
            11'd1110: table_out = 36'hd0b4c9c16;
            11'd1111: table_out = 36'hd0a9956c6;
            11'd1112: table_out = 36'hd09e5ba46;
            11'd1113: table_out = 36'hd0931c644;
            11'd1114: table_out = 36'hd087d7a68;
            11'd1115: table_out = 36'hd07c8d65d;
            11'd1116: table_out = 36'hd0713d9cc;
            11'd1117: table_out = 36'hd065e845f;
            11'd1118: table_out = 36'hd05a8d5bf;
            11'd1119: table_out = 36'hd04f2cd93;
            11'd1120: table_out = 36'hd043c6b82;
            11'd1121: table_out = 36'hd0385af34;
            11'd1122: table_out = 36'hd02ce9850;
            11'd1123: table_out = 36'hd0217267b;
            11'd1124: table_out = 36'hd015f595b;
            11'd1125: table_out = 36'hd00a73095;
            11'd1126: table_out = 36'hcffeeabcd;
            11'd1127: table_out = 36'hcff35caa7;
            11'd1128: table_out = 36'hcfe7c8cc7;
            11'd1129: table_out = 36'hcfdc2f1cf;
            11'd1130: table_out = 36'hcfd08f962;
            11'd1131: table_out = 36'hcfc4ea321;
            11'd1132: table_out = 36'hcfb93eead;
            11'd1133: table_out = 36'hcfad8dba7;
            11'd1134: table_out = 36'hcfa1d69b0;
            11'd1135: table_out = 36'hcf9619865;
            11'd1136: table_out = 36'hcf8a56767;
            11'd1137: table_out = 36'hcf7e8d654;
            11'd1138: table_out = 36'hcf72be4c8;
            11'd1139: table_out = 36'hcf66e9262;
            11'd1140: table_out = 36'hcf5b0debe;
            11'd1141: table_out = 36'hcf4f2c977;
            11'd1142: table_out = 36'hcf434522a;
            11'd1143: table_out = 36'hcf3757870;
            11'd1144: table_out = 36'hcf2b63be4;
            11'd1145: table_out = 36'hcf1f69c1f;
            11'd1146: table_out = 36'hcf13698ba;
            11'd1147: table_out = 36'hcf076314e;
            11'd1148: table_out = 36'hcefb56571;
            11'd1149: table_out = 36'hceef434bb;
            11'd1150: table_out = 36'hcee329ec3;
            11'd1151: table_out = 36'hced70a31d;
            11'd1152: table_out = 36'hcecae415e;
            11'd1153: table_out = 36'hcebeb791c;
            11'd1154: table_out = 36'hceb2849e9;
            11'd1155: table_out = 36'hcea64b358;
            11'd1156: table_out = 36'hce9a0b4fd;
            11'd1157: table_out = 36'hce8dc4e68;
            11'd1158: table_out = 36'hce8177f2a;
            11'd1159: table_out = 36'hce75246d4;
            11'd1160: table_out = 36'hce68ca4f5;
            11'd1161: table_out = 36'hce5c6991c;
            11'd1162: table_out = 36'hce50022d7;
            11'd1163: table_out = 36'hce43941b4;
            11'd1164: table_out = 36'hce371f53f;
            11'd1165: table_out = 36'hce2aa3d03;
            11'd1166: table_out = 36'hce1e2188d;
            11'd1167: table_out = 36'hce1198767;
            11'd1168: table_out = 36'hce050891a;
            11'd1169: table_out = 36'hcdf871d30;
            11'd1170: table_out = 36'hcdebd4330;
            11'd1171: table_out = 36'hcddf2faa1;
            11'd1172: table_out = 36'hcdd28430c;
            11'd1173: table_out = 36'hcdc5d1bf5;
            11'd1174: table_out = 36'hcdb9184e1;
            11'd1175: table_out = 36'hcdac57d55;
            11'd1176: table_out = 36'hcd9f904d5;
            11'd1177: table_out = 36'hcd92c1ae2;
            11'd1178: table_out = 36'hcd85ebeff;
            11'd1179: table_out = 36'hcd790f0ac;
            11'd1180: table_out = 36'hcd6c2af6b;
            11'd1181: table_out = 36'hcd5f3faba;
            11'd1182: table_out = 36'hcd524d218;
            11'd1183: table_out = 36'hcd4553502;
            11'd1184: table_out = 36'hcd38522f5;
            11'd1185: table_out = 36'hcd2b49b6d;
            11'd1186: table_out = 36'hcd1e39de6;
            11'd1187: table_out = 36'hcd11229d9;
            11'd1188: table_out = 36'hcd0403ec0;
            11'd1189: table_out = 36'hccf6ddc12;
            11'd1190: table_out = 36'hcce9b0148;
            11'd1191: table_out = 36'hccdc7add8;
            11'd1192: table_out = 36'hcccf3e138;
            11'd1193: table_out = 36'hccc1f9adc;
            11'd1194: table_out = 36'hccb4ada38;
            11'd1195: table_out = 36'hcca759ebf;
            11'd1196: table_out = 36'hcc99fe7e2;
            11'd1197: table_out = 36'hcc8c9b513;
            11'd1198: table_out = 36'hcc7f305c2;
            11'd1199: table_out = 36'hcc71bd95d;
            11'd1200: table_out = 36'hcc6442f52;
            11'd1201: table_out = 36'hcc56c070f;
            11'd1202: table_out = 36'hcc4935fff;
            11'd1203: table_out = 36'hcc3ba398d;
            11'd1204: table_out = 36'hcc2e09323;
            11'd1205: table_out = 36'hcc2066c29;
            11'd1206: table_out = 36'hcc12bc408;
            11'd1207: table_out = 36'hcc0509a26;
            11'd1208: table_out = 36'hcbf74edea;
            11'd1209: table_out = 36'hcbe98beb6;
            11'd1210: table_out = 36'hcbdbc0bf0;
            11'd1211: table_out = 36'hcbcded4f9;
            11'd1212: table_out = 36'hcbc011933;
            11'd1213: table_out = 36'hcbb22d7fd;
            11'd1214: table_out = 36'hcba4410b7;
            11'd1215: table_out = 36'hcb964c2bf;
            11'd1216: table_out = 36'hcb884ed71;
            11'd1217: table_out = 36'hcb7a49029;
            11'd1218: table_out = 36'hcb6c3aa42;
            11'd1219: table_out = 36'hcb5e23b14;
            11'd1220: table_out = 36'hcb50041f8;
            11'd1221: table_out = 36'hcb41dbe44;
            11'd1222: table_out = 36'hcb33aaf4e;
            11'd1223: table_out = 36'hcb257146b;
            11'd1224: table_out = 36'hcb172eced;
            11'd1225: table_out = 36'hcb08e3826;
            11'd1226: table_out = 36'hcafa8f567;
            11'd1227: table_out = 36'hcaec32400;
            11'd1228: table_out = 36'hcadf26476;
            default : table_out = 36'b0;
        endcase
    end

endmodule