
module inv_shuffle_3 (
    input   [8191:0]  key_shuffle,
    output  [8191:0]  key_original
);
    assign key_original[8191] = key_shuffle[6371];
    assign key_original[8190] = key_shuffle[7935];
    assign key_original[8189] = key_shuffle[5808];
    assign key_original[8188] = key_shuffle[6757];
    assign key_original[8187] = key_shuffle[5659];
    assign key_original[8186] = key_shuffle[6846];
    assign key_original[8185] = key_shuffle[2430];
    assign key_original[8184] = key_shuffle[1816];
    assign key_original[8183] = key_shuffle[3937];
    assign key_original[8182] = key_shuffle[6228];
    assign key_original[8181] = key_shuffle[6273];
    assign key_original[8180] = key_shuffle[4016];
    assign key_original[8179] = key_shuffle[7091];
    assign key_original[8178] = key_shuffle[3555];
    assign key_original[8177] = key_shuffle[4192];
    assign key_original[8176] = key_shuffle[2597];
    assign key_original[8175] = key_shuffle[2079];
    assign key_original[8174] = key_shuffle[6823];
    assign key_original[8173] = key_shuffle[7386];
    assign key_original[8172] = key_shuffle[594];
    assign key_original[8171] = key_shuffle[6359];
    assign key_original[8170] = key_shuffle[7392];
    assign key_original[8169] = key_shuffle[1652];
    assign key_original[8168] = key_shuffle[7335];
    assign key_original[8167] = key_shuffle[4408];
    assign key_original[8166] = key_shuffle[7338];
    assign key_original[8165] = key_shuffle[3803];
    assign key_original[8164] = key_shuffle[4489];
    assign key_original[8163] = key_shuffle[6691];
    assign key_original[8162] = key_shuffle[124];
    assign key_original[8161] = key_shuffle[2725];
    assign key_original[8160] = key_shuffle[2983];
    assign key_original[8159] = key_shuffle[3642];
    assign key_original[8158] = key_shuffle[7944];
    assign key_original[8157] = key_shuffle[7354];
    assign key_original[8156] = key_shuffle[5271];
    assign key_original[8155] = key_shuffle[7771];
    assign key_original[8154] = key_shuffle[3629];
    assign key_original[8153] = key_shuffle[1546];
    assign key_original[8152] = key_shuffle[5047];
    assign key_original[8151] = key_shuffle[570];
    assign key_original[8150] = key_shuffle[5652];
    assign key_original[8149] = key_shuffle[4773];
    assign key_original[8148] = key_shuffle[6424];
    assign key_original[8147] = key_shuffle[4774];
    assign key_original[8146] = key_shuffle[7444];
    assign key_original[8145] = key_shuffle[1047];
    assign key_original[8144] = key_shuffle[5411];
    assign key_original[8143] = key_shuffle[533];
    assign key_original[8142] = key_shuffle[2910];
    assign key_original[8141] = key_shuffle[7680];
    assign key_original[8140] = key_shuffle[4402];
    assign key_original[8139] = key_shuffle[2443];
    assign key_original[8138] = key_shuffle[2619];
    assign key_original[8137] = key_shuffle[7773];
    assign key_original[8136] = key_shuffle[2260];
    assign key_original[8135] = key_shuffle[931];
    assign key_original[8134] = key_shuffle[7941];
    assign key_original[8133] = key_shuffle[1486];
    assign key_original[8132] = key_shuffle[7332];
    assign key_original[8131] = key_shuffle[407];
    assign key_original[8130] = key_shuffle[3256];
    assign key_original[8129] = key_shuffle[3814];
    assign key_original[8128] = key_shuffle[5229];
    assign key_original[8127] = key_shuffle[5821];
    assign key_original[8126] = key_shuffle[5876];
    assign key_original[8125] = key_shuffle[847];
    assign key_original[8124] = key_shuffle[2648];
    assign key_original[8123] = key_shuffle[5549];
    assign key_original[8122] = key_shuffle[7020];
    assign key_original[8121] = key_shuffle[7843];
    assign key_original[8120] = key_shuffle[2627];
    assign key_original[8119] = key_shuffle[6861];
    assign key_original[8118] = key_shuffle[7423];
    assign key_original[8117] = key_shuffle[3026];
    assign key_original[8116] = key_shuffle[7150];
    assign key_original[8115] = key_shuffle[493];
    assign key_original[8114] = key_shuffle[4305];
    assign key_original[8113] = key_shuffle[571];
    assign key_original[8112] = key_shuffle[3796];
    assign key_original[8111] = key_shuffle[3221];
    assign key_original[8110] = key_shuffle[8056];
    assign key_original[8109] = key_shuffle[3299];
    assign key_original[8108] = key_shuffle[1978];
    assign key_original[8107] = key_shuffle[4931];
    assign key_original[8106] = key_shuffle[3064];
    assign key_original[8105] = key_shuffle[5227];
    assign key_original[8104] = key_shuffle[6107];
    assign key_original[8103] = key_shuffle[6601];
    assign key_original[8102] = key_shuffle[4317];
    assign key_original[8101] = key_shuffle[6633];
    assign key_original[8100] = key_shuffle[5507];
    assign key_original[8099] = key_shuffle[6258];
    assign key_original[8098] = key_shuffle[4329];
    assign key_original[8097] = key_shuffle[191];
    assign key_original[8096] = key_shuffle[4002];
    assign key_original[8095] = key_shuffle[1633];
    assign key_original[8094] = key_shuffle[4836];
    assign key_original[8093] = key_shuffle[6738];
    assign key_original[8092] = key_shuffle[2799];
    assign key_original[8091] = key_shuffle[6016];
    assign key_original[8090] = key_shuffle[5011];
    assign key_original[8089] = key_shuffle[2926];
    assign key_original[8088] = key_shuffle[1156];
    assign key_original[8087] = key_shuffle[7654];
    assign key_original[8086] = key_shuffle[1641];
    assign key_original[8085] = key_shuffle[25];
    assign key_original[8084] = key_shuffle[1651];
    assign key_original[8083] = key_shuffle[6151];
    assign key_original[8082] = key_shuffle[4306];
    assign key_original[8081] = key_shuffle[4622];
    assign key_original[8080] = key_shuffle[1438];
    assign key_original[8079] = key_shuffle[6073];
    assign key_original[8078] = key_shuffle[1314];
    assign key_original[8077] = key_shuffle[5823];
    assign key_original[8076] = key_shuffle[953];
    assign key_original[8075] = key_shuffle[1326];
    assign key_original[8074] = key_shuffle[5934];
    assign key_original[8073] = key_shuffle[5314];
    assign key_original[8072] = key_shuffle[3407];
    assign key_original[8071] = key_shuffle[860];
    assign key_original[8070] = key_shuffle[6439];
    assign key_original[8069] = key_shuffle[7696];
    assign key_original[8068] = key_shuffle[6785];
    assign key_original[8067] = key_shuffle[5945];
    assign key_original[8066] = key_shuffle[4001];
    assign key_original[8065] = key_shuffle[6399];
    assign key_original[8064] = key_shuffle[6393];
    assign key_original[8063] = key_shuffle[7699];
    assign key_original[8062] = key_shuffle[147];
    assign key_original[8061] = key_shuffle[730];
    assign key_original[8060] = key_shuffle[3446];
    assign key_original[8059] = key_shuffle[3049];
    assign key_original[8058] = key_shuffle[5706];
    assign key_original[8057] = key_shuffle[2252];
    assign key_original[8056] = key_shuffle[4463];
    assign key_original[8055] = key_shuffle[2241];
    assign key_original[8054] = key_shuffle[6398];
    assign key_original[8053] = key_shuffle[6712];
    assign key_original[8052] = key_shuffle[3747];
    assign key_original[8051] = key_shuffle[1407];
    assign key_original[8050] = key_shuffle[6531];
    assign key_original[8049] = key_shuffle[7263];
    assign key_original[8048] = key_shuffle[6302];
    assign key_original[8047] = key_shuffle[6570];
    assign key_original[8046] = key_shuffle[7714];
    assign key_original[8045] = key_shuffle[1404];
    assign key_original[8044] = key_shuffle[7188];
    assign key_original[8043] = key_shuffle[7130];
    assign key_original[8042] = key_shuffle[1117];
    assign key_original[8041] = key_shuffle[6576];
    assign key_original[8040] = key_shuffle[2809];
    assign key_original[8039] = key_shuffle[6974];
    assign key_original[8038] = key_shuffle[7808];
    assign key_original[8037] = key_shuffle[1479];
    assign key_original[8036] = key_shuffle[2491];
    assign key_original[8035] = key_shuffle[5884];
    assign key_original[8034] = key_shuffle[1799];
    assign key_original[8033] = key_shuffle[6322];
    assign key_original[8032] = key_shuffle[6701];
    assign key_original[8031] = key_shuffle[177];
    assign key_original[8030] = key_shuffle[3176];
    assign key_original[8029] = key_shuffle[7731];
    assign key_original[8028] = key_shuffle[786];
    assign key_original[8027] = key_shuffle[2486];
    assign key_original[8026] = key_shuffle[2483];
    assign key_original[8025] = key_shuffle[1444];
    assign key_original[8024] = key_shuffle[781];
    assign key_original[8023] = key_shuffle[3308];
    assign key_original[8022] = key_shuffle[5729];
    assign key_original[8021] = key_shuffle[5298];
    assign key_original[8020] = key_shuffle[268];
    assign key_original[8019] = key_shuffle[6006];
    assign key_original[8018] = key_shuffle[1756];
    assign key_original[8017] = key_shuffle[7910];
    assign key_original[8016] = key_shuffle[6915];
    assign key_original[8015] = key_shuffle[5971];
    assign key_original[8014] = key_shuffle[2390];
    assign key_original[8013] = key_shuffle[4431];
    assign key_original[8012] = key_shuffle[3916];
    assign key_original[8011] = key_shuffle[3456];
    assign key_original[8010] = key_shuffle[1129];
    assign key_original[8009] = key_shuffle[3263];
    assign key_original[8008] = key_shuffle[3223];
    assign key_original[8007] = key_shuffle[3877];
    assign key_original[8006] = key_shuffle[4838];
    assign key_original[8005] = key_shuffle[5300];
    assign key_original[8004] = key_shuffle[4271];
    assign key_original[8003] = key_shuffle[8103];
    assign key_original[8002] = key_shuffle[7907];
    assign key_original[8001] = key_shuffle[6039];
    assign key_original[8000] = key_shuffle[4521];
    assign key_original[7999] = key_shuffle[5324];
    assign key_original[7998] = key_shuffle[7034];
    assign key_original[7997] = key_shuffle[6419];
    assign key_original[7996] = key_shuffle[7177];
    assign key_original[7995] = key_shuffle[550];
    assign key_original[7994] = key_shuffle[4837];
    assign key_original[7993] = key_shuffle[3587];
    assign key_original[7992] = key_shuffle[7514];
    assign key_original[7991] = key_shuffle[5024];
    assign key_original[7990] = key_shuffle[1913];
    assign key_original[7989] = key_shuffle[6949];
    assign key_original[7988] = key_shuffle[3610];
    assign key_original[7987] = key_shuffle[5294];
    assign key_original[7986] = key_shuffle[254];
    assign key_original[7985] = key_shuffle[3889];
    assign key_original[7984] = key_shuffle[77];
    assign key_original[7983] = key_shuffle[4189];
    assign key_original[7982] = key_shuffle[1053];
    assign key_original[7981] = key_shuffle[6183];
    assign key_original[7980] = key_shuffle[4649];
    assign key_original[7979] = key_shuffle[1764];
    assign key_original[7978] = key_shuffle[6262];
    assign key_original[7977] = key_shuffle[2060];
    assign key_original[7976] = key_shuffle[659];
    assign key_original[7975] = key_shuffle[4602];
    assign key_original[7974] = key_shuffle[4782];
    assign key_original[7973] = key_shuffle[7828];
    assign key_original[7972] = key_shuffle[6810];
    assign key_original[7971] = key_shuffle[6429];
    assign key_original[7970] = key_shuffle[7087];
    assign key_original[7969] = key_shuffle[7809];
    assign key_original[7968] = key_shuffle[881];
    assign key_original[7967] = key_shuffle[5210];
    assign key_original[7966] = key_shuffle[7517];
    assign key_original[7965] = key_shuffle[100];
    assign key_original[7964] = key_shuffle[7649];
    assign key_original[7963] = key_shuffle[4113];
    assign key_original[7962] = key_shuffle[778];
    assign key_original[7961] = key_shuffle[2423];
    assign key_original[7960] = key_shuffle[8168];
    assign key_original[7959] = key_shuffle[2385];
    assign key_original[7958] = key_shuffle[6365];
    assign key_original[7957] = key_shuffle[2520];
    assign key_original[7956] = key_shuffle[3361];
    assign key_original[7955] = key_shuffle[7608];
    assign key_original[7954] = key_shuffle[5514];
    assign key_original[7953] = key_shuffle[7461];
    assign key_original[7952] = key_shuffle[6329];
    assign key_original[7951] = key_shuffle[6580];
    assign key_original[7950] = key_shuffle[2654];
    assign key_original[7949] = key_shuffle[5735];
    assign key_original[7948] = key_shuffle[7549];
    assign key_original[7947] = key_shuffle[3646];
    assign key_original[7946] = key_shuffle[851];
    assign key_original[7945] = key_shuffle[1511];
    assign key_original[7944] = key_shuffle[3312];
    assign key_original[7943] = key_shuffle[2977];
    assign key_original[7942] = key_shuffle[2342];
    assign key_original[7941] = key_shuffle[4904];
    assign key_original[7940] = key_shuffle[3926];
    assign key_original[7939] = key_shuffle[2790];
    assign key_original[7938] = key_shuffle[5822];
    assign key_original[7937] = key_shuffle[3584];
    assign key_original[7936] = key_shuffle[4028];
    assign key_original[7935] = key_shuffle[5569];
    assign key_original[7934] = key_shuffle[7406];
    assign key_original[7933] = key_shuffle[733];
    assign key_original[7932] = key_shuffle[4951];
    assign key_original[7931] = key_shuffle[7664];
    assign key_original[7930] = key_shuffle[3364];
    assign key_original[7929] = key_shuffle[5766];
    assign key_original[7928] = key_shuffle[6314];
    assign key_original[7927] = key_shuffle[3615];
    assign key_original[7926] = key_shuffle[7233];
    assign key_original[7925] = key_shuffle[1239];
    assign key_original[7924] = key_shuffle[4725];
    assign key_original[7923] = key_shuffle[5157];
    assign key_original[7922] = key_shuffle[2287];
    assign key_original[7921] = key_shuffle[4121];
    assign key_original[7920] = key_shuffle[6789];
    assign key_original[7919] = key_shuffle[5562];
    assign key_original[7918] = key_shuffle[6480];
    assign key_original[7917] = key_shuffle[2545];
    assign key_original[7916] = key_shuffle[5343];
    assign key_original[7915] = key_shuffle[7272];
    assign key_original[7914] = key_shuffle[5764];
    assign key_original[7913] = key_shuffle[455];
    assign key_original[7912] = key_shuffle[7298];
    assign key_original[7911] = key_shuffle[704];
    assign key_original[7910] = key_shuffle[1189];
    assign key_original[7909] = key_shuffle[4846];
    assign key_original[7908] = key_shuffle[5902];
    assign key_original[7907] = key_shuffle[2636];
    assign key_original[7906] = key_shuffle[1022];
    assign key_original[7905] = key_shuffle[5690];
    assign key_original[7904] = key_shuffle[1493];
    assign key_original[7903] = key_shuffle[3792];
    assign key_original[7902] = key_shuffle[8021];
    assign key_original[7901] = key_shuffle[5462];
    assign key_original[7900] = key_shuffle[2804];
    assign key_original[7899] = key_shuffle[5548];
    assign key_original[7898] = key_shuffle[5398];
    assign key_original[7897] = key_shuffle[6009];
    assign key_original[7896] = key_shuffle[4719];
    assign key_original[7895] = key_shuffle[4853];
    assign key_original[7894] = key_shuffle[3582];
    assign key_original[7893] = key_shuffle[7072];
    assign key_original[7892] = key_shuffle[6854];
    assign key_original[7891] = key_shuffle[3755];
    assign key_original[7890] = key_shuffle[3295];
    assign key_original[7889] = key_shuffle[639];
    assign key_original[7888] = key_shuffle[899];
    assign key_original[7887] = key_shuffle[8151];
    assign key_original[7886] = key_shuffle[2147];
    assign key_original[7885] = key_shuffle[161];
    assign key_original[7884] = key_shuffle[2614];
    assign key_original[7883] = key_shuffle[7513];
    assign key_original[7882] = key_shuffle[1093];
    assign key_original[7881] = key_shuffle[1952];
    assign key_original[7880] = key_shuffle[6422];
    assign key_original[7879] = key_shuffle[834];
    assign key_original[7878] = key_shuffle[239];
    assign key_original[7877] = key_shuffle[7922];
    assign key_original[7876] = key_shuffle[7747];
    assign key_original[7875] = key_shuffle[2043];
    assign key_original[7874] = key_shuffle[7908];
    assign key_original[7873] = key_shuffle[7707];
    assign key_original[7872] = key_shuffle[5151];
    assign key_original[7871] = key_shuffle[1231];
    assign key_original[7870] = key_shuffle[4675];
    assign key_original[7869] = key_shuffle[2289];
    assign key_original[7868] = key_shuffle[5231];
    assign key_original[7867] = key_shuffle[6857];
    assign key_original[7866] = key_shuffle[4390];
    assign key_original[7865] = key_shuffle[4011];
    assign key_original[7864] = key_shuffle[8128];
    assign key_original[7863] = key_shuffle[2808];
    assign key_original[7862] = key_shuffle[1809];
    assign key_original[7861] = key_shuffle[8026];
    assign key_original[7860] = key_shuffle[6635];
    assign key_original[7859] = key_shuffle[4272];
    assign key_original[7858] = key_shuffle[583];
    assign key_original[7857] = key_shuffle[3258];
    assign key_original[7856] = key_shuffle[4078];
    assign key_original[7855] = key_shuffle[8139];
    assign key_original[7854] = key_shuffle[3536];
    assign key_original[7853] = key_shuffle[5918];
    assign key_original[7852] = key_shuffle[5964];
    assign key_original[7851] = key_shuffle[4713];
    assign key_original[7850] = key_shuffle[1897];
    assign key_original[7849] = key_shuffle[5803];
    assign key_original[7848] = key_shuffle[5956];
    assign key_original[7847] = key_shuffle[5320];
    assign key_original[7846] = key_shuffle[3073];
    assign key_original[7845] = key_shuffle[1869];
    assign key_original[7844] = key_shuffle[8156];
    assign key_original[7843] = key_shuffle[6721];
    assign key_original[7842] = key_shuffle[2153];
    assign key_original[7841] = key_shuffle[5451];
    assign key_original[7840] = key_shuffle[6770];
    assign key_original[7839] = key_shuffle[5740];
    assign key_original[7838] = key_shuffle[8105];
    assign key_original[7837] = key_shuffle[3844];
    assign key_original[7836] = key_shuffle[2444];
    assign key_original[7835] = key_shuffle[7013];
    assign key_original[7834] = key_shuffle[630];
    assign key_original[7833] = key_shuffle[3027];
    assign key_original[7832] = key_shuffle[5301];
    assign key_original[7831] = key_shuffle[43];
    assign key_original[7830] = key_shuffle[377];
    assign key_original[7829] = key_shuffle[7955];
    assign key_original[7828] = key_shuffle[1969];
    assign key_original[7827] = key_shuffle[2204];
    assign key_original[7826] = key_shuffle[1421];
    assign key_original[7825] = key_shuffle[2685];
    assign key_original[7824] = key_shuffle[4917];
    assign key_original[7823] = key_shuffle[3708];
    assign key_original[7822] = key_shuffle[7555];
    assign key_original[7821] = key_shuffle[3112];
    assign key_original[7820] = key_shuffle[2118];
    assign key_original[7819] = key_shuffle[5951];
    assign key_original[7818] = key_shuffle[3124];
    assign key_original[7817] = key_shuffle[4069];
    assign key_original[7816] = key_shuffle[2507];
    assign key_original[7815] = key_shuffle[3502];
    assign key_original[7814] = key_shuffle[4148];
    assign key_original[7813] = key_shuffle[4531];
    assign key_original[7812] = key_shuffle[6549];
    assign key_original[7811] = key_shuffle[2630];
    assign key_original[7810] = key_shuffle[1640];
    assign key_original[7809] = key_shuffle[396];
    assign key_original[7808] = key_shuffle[4099];
    assign key_original[7807] = key_shuffle[1931];
    assign key_original[7806] = key_shuffle[2929];
    assign key_original[7805] = key_shuffle[7044];
    assign key_original[7804] = key_shuffle[1051];
    assign key_original[7803] = key_shuffle[6684];
    assign key_original[7802] = key_shuffle[2684];
    assign key_original[7801] = key_shuffle[4278];
    assign key_original[7800] = key_shuffle[3857];
    assign key_original[7799] = key_shuffle[7848];
    assign key_original[7798] = key_shuffle[1337];
    assign key_original[7797] = key_shuffle[1149];
    assign key_original[7796] = key_shuffle[1745];
    assign key_original[7795] = key_shuffle[5388];
    assign key_original[7794] = key_shuffle[4426];
    assign key_original[7793] = key_shuffle[1808];
    assign key_original[7792] = key_shuffle[2398];
    assign key_original[7791] = key_shuffle[266];
    assign key_original[7790] = key_shuffle[1776];
    assign key_original[7789] = key_shuffle[5495];
    assign key_original[7788] = key_shuffle[5027];
    assign key_original[7787] = key_shuffle[3975];
    assign key_original[7786] = key_shuffle[6535];
    assign key_original[7785] = key_shuffle[7510];
    assign key_original[7784] = key_shuffle[7830];
    assign key_original[7783] = key_shuffle[4549];
    assign key_original[7782] = key_shuffle[6323];
    assign key_original[7781] = key_shuffle[6594];
    assign key_original[7780] = key_shuffle[6603];
    assign key_original[7779] = key_shuffle[3097];
    assign key_original[7778] = key_shuffle[993];
    assign key_original[7777] = key_shuffle[5353];
    assign key_original[7776] = key_shuffle[4486];
    assign key_original[7775] = key_shuffle[4687];
    assign key_original[7774] = key_shuffle[5637];
    assign key_original[7773] = key_shuffle[6845];
    assign key_original[7772] = key_shuffle[891];
    assign key_original[7771] = key_shuffle[419];
    assign key_original[7770] = key_shuffle[8114];
    assign key_original[7769] = key_shuffle[3437];
    assign key_original[7768] = key_shuffle[4356];
    assign key_original[7767] = key_shuffle[5241];
    assign key_original[7766] = key_shuffle[1713];
    assign key_original[7765] = key_shuffle[6078];
    assign key_original[7764] = key_shuffle[1695];
    assign key_original[7763] = key_shuffle[295];
    assign key_original[7762] = key_shuffle[90];
    assign key_original[7761] = key_shuffle[272];
    assign key_original[7760] = key_shuffle[5268];
    assign key_original[7759] = key_shuffle[6578];
    assign key_original[7758] = key_shuffle[912];
    assign key_original[7757] = key_shuffle[1797];
    assign key_original[7756] = key_shuffle[6912];
    assign key_original[7755] = key_shuffle[5614];
    assign key_original[7754] = key_shuffle[1852];
    assign key_original[7753] = key_shuffle[3072];
    assign key_original[7752] = key_shuffle[2884];
    assign key_original[7751] = key_shuffle[2127];
    assign key_original[7750] = key_shuffle[3215];
    assign key_original[7749] = key_shuffle[3746];
    assign key_original[7748] = key_shuffle[6819];
    assign key_original[7747] = key_shuffle[7739];
    assign key_original[7746] = key_shuffle[517];
    assign key_original[7745] = key_shuffle[7964];
    assign key_original[7744] = key_shuffle[6119];
    assign key_original[7743] = key_shuffle[5634];
    assign key_original[7742] = key_shuffle[4047];
    assign key_original[7741] = key_shuffle[3578];
    assign key_original[7740] = key_shuffle[5051];
    assign key_original[7739] = key_shuffle[6376];
    assign key_original[7738] = key_shuffle[2975];
    assign key_original[7737] = key_shuffle[3421];
    assign key_original[7736] = key_shuffle[880];
    assign key_original[7735] = key_shuffle[2878];
    assign key_original[7734] = key_shuffle[3621];
    assign key_original[7733] = key_shuffle[6938];
    assign key_original[7732] = key_shuffle[1161];
    assign key_original[7731] = key_shuffle[6847];
    assign key_original[7730] = key_shuffle[6648];
    assign key_original[7729] = key_shuffle[7080];
    assign key_original[7728] = key_shuffle[6650];
    assign key_original[7727] = key_shuffle[5250];
    assign key_original[7726] = key_shuffle[747];
    assign key_original[7725] = key_shuffle[4615];
    assign key_original[7724] = key_shuffle[4511];
    assign key_original[7723] = key_shuffle[1204];
    assign key_original[7722] = key_shuffle[2886];
    assign key_original[7721] = key_shuffle[6844];
    assign key_original[7720] = key_shuffle[3870];
    assign key_original[7719] = key_shuffle[5248];
    assign key_original[7718] = key_shuffle[4216];
    assign key_original[7717] = key_shuffle[4660];
    assign key_original[7716] = key_shuffle[1953];
    assign key_original[7715] = key_shuffle[703];
    assign key_original[7714] = key_shuffle[7028];
    assign key_original[7713] = key_shuffle[3867];
    assign key_original[7712] = key_shuffle[6289];
    assign key_original[7711] = key_shuffle[7276];
    assign key_original[7710] = key_shuffle[3423];
    assign key_original[7709] = key_shuffle[5194];
    assign key_original[7708] = key_shuffle[6715];
    assign key_original[7707] = key_shuffle[6920];
    assign key_original[7706] = key_shuffle[4409];
    assign key_original[7705] = key_shuffle[4810];
    assign key_original[7704] = key_shuffle[4668];
    assign key_original[7703] = key_shuffle[753];
    assign key_original[7702] = key_shuffle[7221];
    assign key_original[7701] = key_shuffle[7388];
    assign key_original[7700] = key_shuffle[6063];
    assign key_original[7699] = key_shuffle[2776];
    assign key_original[7698] = key_shuffle[60];
    assign key_original[7697] = key_shuffle[3368];
    assign key_original[7696] = key_shuffle[845];
    assign key_original[7695] = key_shuffle[2535];
    assign key_original[7694] = key_shuffle[1375];
    assign key_original[7693] = key_shuffle[4913];
    assign key_original[7692] = key_shuffle[4624];
    assign key_original[7691] = key_shuffle[600];
    assign key_original[7690] = key_shuffle[3428];
    assign key_original[7689] = key_shuffle[7596];
    assign key_original[7688] = key_shuffle[7323];
    assign key_original[7687] = key_shuffle[3560];
    assign key_original[7686] = key_shuffle[898];
    assign key_original[7685] = key_shuffle[6379];
    assign key_original[7684] = key_shuffle[3068];
    assign key_original[7683] = key_shuffle[5708];
    assign key_original[7682] = key_shuffle[1387];
    assign key_original[7681] = key_shuffle[3400];
    assign key_original[7680] = key_shuffle[3509];
    assign key_original[7679] = key_shuffle[3189];
    assign key_original[7678] = key_shuffle[6342];
    assign key_original[7677] = key_shuffle[8174];
    assign key_original[7676] = key_shuffle[1446];
    assign key_original[7675] = key_shuffle[3960];
    assign key_original[7674] = key_shuffle[6527];
    assign key_original[7673] = key_shuffle[1624];
    assign key_original[7672] = key_shuffle[5376];
    assign key_original[7671] = key_shuffle[2540];
    assign key_original[7670] = key_shuffle[1440];
    assign key_original[7669] = key_shuffle[7946];
    assign key_original[7668] = key_shuffle[5895];
    assign key_original[7667] = key_shuffle[6361];
    assign key_original[7666] = key_shuffle[6795];
    assign key_original[7665] = key_shuffle[7264];
    assign key_original[7664] = key_shuffle[940];
    assign key_original[7663] = key_shuffle[1081];
    assign key_original[7662] = key_shuffle[4753];
    assign key_original[7661] = key_shuffle[2005];
    assign key_original[7660] = key_shuffle[7404];
    assign key_original[7659] = key_shuffle[863];
    assign key_original[7658] = key_shuffle[3904];
    assign key_original[7657] = key_shuffle[1233];
    assign key_original[7656] = key_shuffle[6799];
    assign key_original[7655] = key_shuffle[6689];
    assign key_original[7654] = key_shuffle[5969];
    assign key_original[7653] = key_shuffle[5568];
    assign key_original[7652] = key_shuffle[7101];
    assign key_original[7651] = key_shuffle[5463];
    assign key_original[7650] = key_shuffle[3931];
    assign key_original[7649] = key_shuffle[3067];
    assign key_original[7648] = key_shuffle[5312];
    assign key_original[7647] = key_shuffle[6654];
    assign key_original[7646] = key_shuffle[12];
    assign key_original[7645] = key_shuffle[2090];
    assign key_original[7644] = key_shuffle[5788];
    assign key_original[7643] = key_shuffle[4459];
    assign key_original[7642] = key_shuffle[1418];
    assign key_original[7641] = key_shuffle[5050];
    assign key_original[7640] = key_shuffle[3012];
    assign key_original[7639] = key_shuffle[1230];
    assign key_original[7638] = key_shuffle[5838];
    assign key_original[7637] = key_shuffle[5641];
    assign key_original[7636] = key_shuffle[4737];
    assign key_original[7635] = key_shuffle[3199];
    assign key_original[7634] = key_shuffle[7879];
    assign key_original[7633] = key_shuffle[243];
    assign key_original[7632] = key_shuffle[4590];
    assign key_original[7631] = key_shuffle[8167];
    assign key_original[7630] = key_shuffle[5391];
    assign key_original[7629] = key_shuffle[3138];
    assign key_original[7628] = key_shuffle[2850];
    assign key_original[7627] = key_shuffle[6478];
    assign key_original[7626] = key_shuffle[929];
    assign key_original[7625] = key_shuffle[5778];
    assign key_original[7624] = key_shuffle[8054];
    assign key_original[7623] = key_shuffle[2816];
    assign key_original[7622] = key_shuffle[7791];
    assign key_original[7621] = key_shuffle[5371];
    assign key_original[7620] = key_shuffle[652];
    assign key_original[7619] = key_shuffle[5364];
    assign key_original[7618] = key_shuffle[3195];
    assign key_original[7617] = key_shuffle[6908];
    assign key_original[7616] = key_shuffle[4971];
    assign key_original[7615] = key_shuffle[1674];
    assign key_original[7614] = key_shuffle[6832];
    assign key_original[7613] = key_shuffle[4674];
    assign key_original[7612] = key_shuffle[1172];
    assign key_original[7611] = key_shuffle[7966];
    assign key_original[7610] = key_shuffle[7496];
    assign key_original[7609] = key_shuffle[4678];
    assign key_original[7608] = key_shuffle[7711];
    assign key_original[7607] = key_shuffle[4088];
    assign key_original[7606] = key_shuffle[3962];
    assign key_original[7605] = key_shuffle[8033];
    assign key_original[7604] = key_shuffle[1773];
    assign key_original[7603] = key_shuffle[2462];
    assign key_original[7602] = key_shuffle[1174];
    assign key_original[7601] = key_shuffle[333];
    assign key_original[7600] = key_shuffle[7036];
    assign key_original[7599] = key_shuffle[3153];
    assign key_original[7598] = key_shuffle[815];
    assign key_original[7597] = key_shuffle[7916];
    assign key_original[7596] = key_shuffle[2557];
    assign key_original[7595] = key_shuffle[1202];
    assign key_original[7594] = key_shuffle[6867];
    assign key_original[7593] = key_shuffle[2202];
    assign key_original[7592] = key_shuffle[1247];
    assign key_original[7591] = key_shuffle[1775];
    assign key_original[7590] = key_shuffle[1428];
    assign key_original[7589] = key_shuffle[5503];
    assign key_original[7588] = key_shuffle[6952];
    assign key_original[7587] = key_shuffle[5406];
    assign key_original[7586] = key_shuffle[2938];
    assign key_original[7585] = key_shuffle[5912];
    assign key_original[7584] = key_shuffle[6640];
    assign key_original[7583] = key_shuffle[7862];
    assign key_original[7582] = key_shuffle[3283];
    assign key_original[7581] = key_shuffle[1103];
    assign key_original[7580] = key_shuffle[4518];
    assign key_original[7579] = key_shuffle[4095];
    assign key_original[7578] = key_shuffle[769];
    assign key_original[7577] = key_shuffle[2715];
    assign key_original[7576] = key_shuffle[2242];
    assign key_original[7575] = key_shuffle[1538];
    assign key_original[7574] = key_shuffle[4140];
    assign key_original[7573] = key_shuffle[6448];
    assign key_original[7572] = key_shuffle[6541];
    assign key_original[7571] = key_shuffle[3311];
    assign key_original[7570] = key_shuffle[4224];
    assign key_original[7569] = key_shuffle[4962];
    assign key_original[7568] = key_shuffle[660];
    assign key_original[7567] = key_shuffle[6416];
    assign key_original[7566] = key_shuffle[7833];
    assign key_original[7565] = key_shuffle[3110];
    assign key_original[7564] = key_shuffle[143];
    assign key_original[7563] = key_shuffle[1561];
    assign key_original[7562] = key_shuffle[7651];
    assign key_original[7561] = key_shuffle[4249];
    assign key_original[7560] = key_shuffle[2472];
    assign key_original[7559] = key_shuffle[6030];
    assign key_original[7558] = key_shuffle[5703];
    assign key_original[7557] = key_shuffle[2963];
    assign key_original[7556] = key_shuffle[6765];
    assign key_original[7555] = key_shuffle[1787];
    assign key_original[7554] = key_shuffle[5830];
    assign key_original[7553] = key_shuffle[2839];
    assign key_original[7552] = key_shuffle[5714];
    assign key_original[7551] = key_shuffle[2997];
    assign key_original[7550] = key_shuffle[5362];
    assign key_original[7549] = key_shuffle[3147];
    assign key_original[7548] = key_shuffle[1448];
    assign key_original[7547] = key_shuffle[889];
    assign key_original[7546] = key_shuffle[2500];
    assign key_original[7545] = key_shuffle[5150];
    assign key_original[7544] = key_shuffle[3477];
    assign key_original[7543] = key_shuffle[1499];
    assign key_original[7542] = key_shuffle[8140];
    assign key_original[7541] = key_shuffle[7352];
    assign key_original[7540] = key_shuffle[2180];
    assign key_original[7539] = key_shuffle[2524];
    assign key_original[7538] = key_shuffle[4763];
    assign key_original[7537] = key_shuffle[4591];
    assign key_original[7536] = key_shuffle[3066];
    assign key_original[7535] = key_shuffle[2115];
    assign key_original[7534] = key_shuffle[3057];
    assign key_original[7533] = key_shuffle[2814];
    assign key_original[7532] = key_shuffle[74];
    assign key_original[7531] = key_shuffle[7210];
    assign key_original[7530] = key_shuffle[47];
    assign key_original[7529] = key_shuffle[3710];
    assign key_original[7528] = key_shuffle[5925];
    assign key_original[7527] = key_shuffle[1323];
    assign key_original[7526] = key_shuffle[1414];
    assign key_original[7525] = key_shuffle[3725];
    assign key_original[7524] = key_shuffle[2463];
    assign key_original[7523] = key_shuffle[6112];
    assign key_original[7522] = key_shuffle[8191];
    assign key_original[7521] = key_shuffle[5528];
    assign key_original[7520] = key_shuffle[7222];
    assign key_original[7519] = key_shuffle[3166];
    assign key_original[7518] = key_shuffle[5267];
    assign key_original[7517] = key_shuffle[4950];
    assign key_original[7516] = key_shuffle[2730];
    assign key_original[7515] = key_shuffle[6997];
    assign key_original[7514] = key_shuffle[4808];
    assign key_original[7513] = key_shuffle[3322];
    assign key_original[7512] = key_shuffle[3512];
    assign key_original[7511] = key_shuffle[6042];
    assign key_original[7510] = key_shuffle[2410];
    assign key_original[7509] = key_shuffle[1220];
    assign key_original[7508] = key_shuffle[7416];
    assign key_original[7507] = key_shuffle[866];
    assign key_original[7506] = key_shuffle[1580];
    assign key_original[7505] = key_shuffle[7566];
    assign key_original[7504] = key_shuffle[1662];
    assign key_original[7503] = key_shuffle[5214];
    assign key_original[7502] = key_shuffle[8089];
    assign key_original[7501] = key_shuffle[710];
    assign key_original[7500] = key_shuffle[6816];
    assign key_original[7499] = key_shuffle[6315];
    assign key_original[7498] = key_shuffle[2341];
    assign key_original[7497] = key_shuffle[7076];
    assign key_original[7496] = key_shuffle[3109];
    assign key_original[7495] = key_shuffle[7390];
    assign key_original[7494] = key_shuffle[873];
    assign key_original[7493] = key_shuffle[4710];
    assign key_original[7492] = key_shuffle[7567];
    assign key_original[7491] = key_shuffle[69];
    assign key_original[7490] = key_shuffle[2259];
    assign key_original[7489] = key_shuffle[3020];
    assign key_original[7488] = key_shuffle[2643];
    assign key_original[7487] = key_shuffle[5663];
    assign key_original[7486] = key_shuffle[5017];
    assign key_original[7485] = key_shuffle[6951];
    assign key_original[7484] = key_shuffle[6564];
    assign key_original[7483] = key_shuffle[5741];
    assign key_original[7482] = key_shuffle[5639];
    assign key_original[7481] = key_shuffle[6887];
    assign key_original[7480] = key_shuffle[1134];
    assign key_original[7479] = key_shuffle[4446];
    assign key_original[7478] = key_shuffle[7421];
    assign key_original[7477] = key_shuffle[4132];
    assign key_original[7476] = key_shuffle[745];
    assign key_original[7475] = key_shuffle[6970];
    assign key_original[7474] = key_shuffle[4115];
    assign key_original[7473] = key_shuffle[5344];
    assign key_original[7472] = key_shuffle[8148];
    assign key_original[7471] = key_shuffle[8001];
    assign key_original[7470] = key_shuffle[1271];
    assign key_original[7469] = key_shuffle[3565];
    assign key_original[7468] = key_shuffle[4371];
    assign key_original[7467] = key_shuffle[7112];
    assign key_original[7466] = key_shuffle[1955];
    assign key_original[7465] = key_shuffle[1012];
    assign key_original[7464] = key_shuffle[3301];
    assign key_original[7463] = key_shuffle[4625];
    assign key_original[7462] = key_shuffle[3817];
    assign key_original[7461] = key_shuffle[4400];
    assign key_original[7460] = key_shuffle[1069];
    assign key_original[7459] = key_shuffle[2250];
    assign key_original[7458] = key_shuffle[6412];
    assign key_original[7457] = key_shuffle[5588];
    assign key_original[7456] = key_shuffle[1579];
    assign key_original[7455] = key_shuffle[53];
    assign key_original[7454] = key_shuffle[87];
    assign key_original[7453] = key_shuffle[7986];
    assign key_original[7452] = key_shuffle[982];
    assign key_original[7451] = key_shuffle[2902];
    assign key_original[7450] = key_shuffle[2510];
    assign key_original[7449] = key_shuffle[5733];
    assign key_original[7448] = key_shuffle[417];
    assign key_original[7447] = key_shuffle[6259];
    assign key_original[7446] = key_shuffle[6745];
    assign key_original[7445] = key_shuffle[4474];
    assign key_original[7444] = key_shuffle[3805];
    assign key_original[7443] = key_shuffle[7448];
    assign key_original[7442] = key_shuffle[1263];
    assign key_original[7441] = key_shuffle[6964];
    assign key_original[7440] = key_shuffle[6240];
    assign key_original[7439] = key_shuffle[6822];
    assign key_original[7438] = key_shuffle[7762];
    assign key_original[7437] = key_shuffle[1360];
    assign key_original[7436] = key_shuffle[1549];
    assign key_original[7435] = key_shuffle[2040];
    assign key_original[7434] = key_shuffle[2863];
    assign key_original[7433] = key_shuffle[4857];
    assign key_original[7432] = key_shuffle[7719];
    assign key_original[7431] = key_shuffle[349];
    assign key_original[7430] = key_shuffle[2205];
    assign key_original[7429] = key_shuffle[7744];
    assign key_original[7428] = key_shuffle[7702];
    assign key_original[7427] = key_shuffle[4886];
    assign key_original[7426] = key_shuffle[155];
    assign key_original[7425] = key_shuffle[2309];
    assign key_original[7424] = key_shuffle[224];
    assign key_original[7423] = key_shuffle[4733];
    assign key_original[7422] = key_shuffle[2968];
    assign key_original[7421] = key_shuffle[7413];
    assign key_original[7420] = key_shuffle[6307];
    assign key_original[7419] = key_shuffle[5923];
    assign key_original[7418] = key_shuffle[638];
    assign key_original[7417] = key_shuffle[2571];
    assign key_original[7416] = key_shuffle[3239];
    assign key_original[7415] = key_shuffle[4363];
    assign key_original[7414] = key_shuffle[6708];
    assign key_original[7413] = key_shuffle[7086];
    assign key_original[7412] = key_shuffle[7898];
    assign key_original[7411] = key_shuffle[6346];
    assign key_original[7410] = key_shuffle[6265];
    assign key_original[7409] = key_shuffle[3516];
    assign key_original[7408] = key_shuffle[3680];
    assign key_original[7407] = key_shuffle[2862];
    assign key_original[7406] = key_shuffle[6225];
    assign key_original[7405] = key_shuffle[6312];
    assign key_original[7404] = key_shuffle[1827];
    assign key_original[7403] = key_shuffle[7793];
    assign key_original[7402] = key_shuffle[1982];
    assign key_original[7401] = key_shuffle[7228];
    assign key_original[7400] = key_shuffle[4706];
    assign key_original[7399] = key_shuffle[4333];
    assign key_original[7398] = key_shuffle[1628];
    assign key_original[7397] = key_shuffle[7303];
    assign key_original[7396] = key_shuffle[7743];
    assign key_original[7395] = key_shuffle[1339];
    assign key_original[7394] = key_shuffle[4750];
    assign key_original[7393] = key_shuffle[3608];
    assign key_original[7392] = key_shuffle[492];
    assign key_original[7391] = key_shuffle[6537];
    assign key_original[7390] = key_shuffle[5474];
    assign key_original[7389] = key_shuffle[4199];
    assign key_original[7388] = key_shuffle[3129];
    assign key_original[7387] = key_shuffle[7414];
    assign key_original[7386] = key_shuffle[1291];
    assign key_original[7385] = key_shuffle[1926];
    assign key_original[7384] = key_shuffle[6066];
    assign key_original[7383] = key_shuffle[4947];
    assign key_original[7382] = key_shuffle[2930];
    assign key_original[7381] = key_shuffle[4049];
    assign key_original[7380] = key_shuffle[4514];
    assign key_original[7379] = key_shuffle[1322];
    assign key_original[7378] = key_shuffle[7271];
    assign key_original[7377] = key_shuffle[1536];
    assign key_original[7376] = key_shuffle[1473];
    assign key_original[7375] = key_shuffle[5797];
    assign key_original[7374] = key_shuffle[1942];
    assign key_original[7373] = key_shuffle[5942];
    assign key_original[7372] = key_shuffle[817];
    assign key_original[7371] = key_shuffle[5546];
    assign key_original[7370] = key_shuffle[540];
    assign key_original[7369] = key_shuffle[5502];
    assign key_original[7368] = key_shuffle[1253];
    assign key_original[7367] = key_shuffle[4863];
    assign key_original[7366] = key_shuffle[1627];
    assign key_original[7365] = key_shuffle[5119];
    assign key_original[7364] = key_shuffle[6291];
    assign key_original[7363] = key_shuffle[6807];
    assign key_original[7362] = key_shuffle[7174];
    assign key_original[7361] = key_shuffle[2695];
    assign key_original[7360] = key_shuffle[2015];
    assign key_original[7359] = key_shuffle[1201];
    assign key_original[7358] = key_shuffle[5366];
    assign key_original[7357] = key_shuffle[4623];
    assign key_original[7356] = key_shuffle[6522];
    assign key_original[7355] = key_shuffle[6797];
    assign key_original[7354] = key_shuffle[8189];
    assign key_original[7353] = key_shuffle[5083];
    assign key_original[7352] = key_shuffle[4039];
    assign key_original[7351] = key_shuffle[4898];
    assign key_original[7350] = key_shuffle[8127];
    assign key_original[7349] = key_shuffle[237];
    assign key_original[7348] = key_shuffle[7796];
    assign key_original[7347] = key_shuffle[1551];
    assign key_original[7346] = key_shuffle[910];
    assign key_original[7345] = key_shuffle[5532];
    assign key_original[7344] = key_shuffle[6834];
    assign key_original[7343] = key_shuffle[3077];
    assign key_original[7342] = key_shuffle[1564];
    assign key_original[7341] = key_shuffle[1282];
    assign key_original[7340] = key_shuffle[6029];
    assign key_original[7339] = key_shuffle[4594];
    assign key_original[7338] = key_shuffle[7780];
    assign key_original[7337] = key_shuffle[1613];
    assign key_original[7336] = key_shuffle[8099];
    assign key_original[7335] = key_shuffle[7190];
    assign key_original[7334] = key_shuffle[11];
    assign key_original[7333] = key_shuffle[7176];
    assign key_original[7332] = key_shuffle[3469];
    assign key_original[7331] = key_shuffle[7670];
    assign key_original[7330] = key_shuffle[5579];
    assign key_original[7329] = key_shuffle[2859];
    assign key_original[7328] = key_shuffle[7669];
    assign key_original[7327] = key_shuffle[7952];
    assign key_original[7326] = key_shuffle[1084];
    assign key_original[7325] = key_shuffle[5232];
    assign key_original[7324] = key_shuffle[5352];
    assign key_original[7323] = key_shuffle[7327];
    assign key_original[7322] = key_shuffle[7724];
    assign key_original[7321] = key_shuffle[3942];
    assign key_original[7320] = key_shuffle[7591];
    assign key_original[7319] = key_shuffle[3993];
    assign key_original[7318] = key_shuffle[6319];
    assign key_original[7317] = key_shuffle[2251];
    assign key_original[7316] = key_shuffle[4676];
    assign key_original[7315] = key_shuffle[2319];
    assign key_original[7314] = key_shuffle[2948];
    assign key_original[7313] = key_shuffle[3598];
    assign key_original[7312] = key_shuffle[1324];
    assign key_original[7311] = key_shuffle[4578];
    assign key_original[7310] = key_shuffle[7900];
    assign key_original[7309] = key_shuffle[3000];
    assign key_original[7308] = key_shuffle[556];
    assign key_original[7307] = key_shuffle[4480];
    assign key_original[7306] = key_shuffle[3174];
    assign key_original[7305] = key_shuffle[6994];
    assign key_original[7304] = key_shuffle[3201];
    assign key_original[7303] = key_shuffle[5221];
    assign key_original[7302] = key_shuffle[2517];
    assign key_original[7301] = key_shuffle[4819];
    assign key_original[7300] = key_shuffle[7074];
    assign key_original[7299] = key_shuffle[3932];
    assign key_original[7298] = key_shuffle[890];
    assign key_original[7297] = key_shuffle[7522];
    assign key_original[7296] = key_shuffle[1240];
    assign key_original[7295] = key_shuffle[2460];
    assign key_original[7294] = key_shuffle[3481];
    assign key_original[7293] = key_shuffle[3045];
    assign key_original[7292] = key_shuffle[7620];
    assign key_original[7291] = key_shuffle[7380];
    assign key_original[7290] = key_shuffle[3611];
    assign key_original[7289] = key_shuffle[2602];
    assign key_original[7288] = key_shuffle[821];
    assign key_original[7287] = key_shuffle[8117];
    assign key_original[7286] = key_shuffle[5377];
    assign key_original[7285] = key_shuffle[4154];
    assign key_original[7284] = key_shuffle[2455];
    assign key_original[7283] = key_shuffle[3620];
    assign key_original[7282] = key_shuffle[8022];
    assign key_original[7281] = key_shuffle[542];
    assign key_original[7280] = key_shuffle[7798];
    assign key_original[7279] = key_shuffle[7218];
    assign key_original[7278] = key_shuffle[3868];
    assign key_original[7277] = key_shuffle[6750];
    assign key_original[7276] = key_shuffle[2349];
    assign key_original[7275] = key_shuffle[4484];
    assign key_original[7274] = key_shuffle[2206];
    assign key_original[7273] = key_shuffle[666];
    assign key_original[7272] = key_shuffle[2758];
    assign key_original[7271] = key_shuffle[133];
    assign key_original[7270] = key_shuffle[379];
    assign key_original[7269] = key_shuffle[7580];
    assign key_original[7268] = key_shuffle[4876];
    assign key_original[7267] = key_shuffle[2764];
    assign key_original[7266] = key_shuffle[6249];
    assign key_original[7265] = key_shuffle[6100];
    assign key_original[7264] = key_shuffle[5787];
    assign key_original[7263] = key_shuffle[2606];
    assign key_original[7262] = key_shuffle[5886];
    assign key_original[7261] = key_shuffle[1672];
    assign key_original[7260] = key_shuffle[1772];
    assign key_original[7259] = key_shuffle[6226];
    assign key_original[7258] = key_shuffle[2547];
    assign key_original[7257] = key_shuffle[987];
    assign key_original[7256] = key_shuffle[1987];
    assign key_original[7255] = key_shuffle[4924];
    assign key_original[7254] = key_shuffle[317];
    assign key_original[7253] = key_shuffle[1889];
    assign key_original[7252] = key_shuffle[7260];
    assign key_original[7251] = key_shuffle[3168];
    assign key_original[7250] = key_shuffle[2513];
    assign key_original[7249] = key_shuffle[838];
    assign key_original[7248] = key_shuffle[7979];
    assign key_original[7247] = key_shuffle[3396];
    assign key_original[7246] = key_shuffle[1607];
    assign key_original[7245] = key_shuffle[2176];
    assign key_original[7244] = key_shuffle[1487];
    assign key_original[7243] = key_shuffle[5443];
    assign key_original[7242] = key_shuffle[6043];
    assign key_original[7241] = key_shuffle[2297];
    assign key_original[7240] = key_shuffle[5916];
    assign key_original[7239] = key_shuffle[6054];
    assign key_original[7238] = key_shuffle[7313];
    assign key_original[7237] = key_shuffle[1210];
    assign key_original[7236] = key_shuffle[6058];
    assign key_original[7235] = key_shuffle[2021];
    assign key_original[7234] = key_shuffle[4646];
    assign key_original[7233] = key_shuffle[7838];
    assign key_original[7232] = key_shuffle[5878];
    assign key_original[7231] = key_shuffle[4565];
    assign key_original[7230] = key_shuffle[2953];
    assign key_original[7229] = key_shuffle[2693];
    assign key_original[7228] = key_shuffle[5274];
    assign key_original[7227] = key_shuffle[4157];
    assign key_original[7226] = key_shuffle[1752];
    assign key_original[7225] = key_shuffle[7379];
    assign key_original[7224] = key_shuffle[8053];
    assign key_original[7223] = key_shuffle[7950];
    assign key_original[7222] = key_shuffle[4516];
    assign key_original[7221] = key_shuffle[4970];
    assign key_original[7220] = key_shuffle[6598];
    assign key_original[7219] = key_shuffle[3131];
    assign key_original[7218] = key_shuffle[4783];
    assign key_original[7217] = key_shuffle[1941];
    assign key_original[7216] = key_shuffle[1112];
    assign key_original[7215] = key_shuffle[390];
    assign key_original[7214] = key_shuffle[7867];
    assign key_original[7213] = key_shuffle[5561];
    assign key_original[7212] = key_shuffle[7643];
    assign key_original[7211] = key_shuffle[5422];
    assign key_original[7210] = key_shuffle[4659];
    assign key_original[7209] = key_shuffle[3259];
    assign key_original[7208] = key_shuffle[4070];
    assign key_original[7207] = key_shuffle[180];
    assign key_original[7206] = key_shuffle[3544];
    assign key_original[7205] = key_shuffle[4989];
    assign key_original[7204] = key_shuffle[530];
    assign key_original[7203] = key_shuffle[3827];
    assign key_original[7202] = key_shuffle[5727];
    assign key_original[7201] = key_shuffle[2171];
    assign key_original[7200] = key_shuffle[4688];
    assign key_original[7199] = key_shuffle[6162];
    assign key_original[7198] = key_shuffle[6330];
    assign key_original[7197] = key_shuffle[2958];
    assign key_original[7196] = key_shuffle[3466];
    assign key_original[7195] = key_shuffle[3525];
    assign key_original[7194] = key_shuffle[356];
    assign key_original[7193] = key_shuffle[4059];
    assign key_original[7192] = key_shuffle[7903];
    assign key_original[7191] = key_shuffle[7556];
    assign key_original[7190] = key_shuffle[4546];
    assign key_original[7189] = key_shuffle[1005];
    assign key_original[7188] = key_shuffle[5078];
    assign key_original[7187] = key_shuffle[2563];
    assign key_original[7186] = key_shuffle[3531];
    assign key_original[7185] = key_shuffle[4842];
    assign key_original[7184] = key_shuffle[2312];
    assign key_original[7183] = key_shuffle[7241];
    assign key_original[7182] = key_shuffle[4419];
    assign key_original[7181] = key_shuffle[6793];
    assign key_original[7180] = key_shuffle[8078];
    assign key_original[7179] = key_shuffle[3595];
    assign key_original[7178] = key_shuffle[7569];
    assign key_original[7177] = key_shuffle[1895];
    assign key_original[7176] = key_shuffle[3949];
    assign key_original[7175] = key_shuffle[4526];
    assign key_original[7174] = key_shuffle[687];
    assign key_original[7173] = key_shuffle[6554];
    assign key_original[7172] = key_shuffle[2689];
    assign key_original[7171] = key_shuffle[5527];
    assign key_original[7170] = key_shuffle[7752];
    assign key_original[7169] = key_shuffle[6548];
    assign key_original[7168] = key_shuffle[5099];
    assign key_original[7167] = key_shuffle[136];
    assign key_original[7166] = key_shuffle[3718];
    assign key_original[7165] = key_shuffle[7819];
    assign key_original[7164] = key_shuffle[3639];
    assign key_original[7163] = key_shuffle[598];
    assign key_original[7162] = key_shuffle[4455];
    assign key_original[7161] = key_shuffle[2714];
    assign key_original[7160] = key_shuffle[3117];
    assign key_original[7159] = key_shuffle[5147];
    assign key_original[7158] = key_shuffle[3722];
    assign key_original[7157] = key_shuffle[2591];
    assign key_original[7156] = key_shuffle[4407];
    assign key_original[7155] = key_shuffle[1635];
    assign key_original[7154] = key_shuffle[7251];
    assign key_original[7153] = key_shuffle[5691];
    assign key_original[7152] = key_shuffle[5068];
    assign key_original[7151] = key_shuffle[3211];
    assign key_original[7150] = key_shuffle[4227];
    assign key_original[7149] = key_shuffle[4722];
    assign key_original[7148] = key_shuffle[3963];
    assign key_original[7147] = key_shuffle[3365];
    assign key_original[7146] = key_shuffle[1075];
    assign key_original[7145] = key_shuffle[5784];
    assign key_original[7144] = key_shuffle[1356];
    assign key_original[7143] = key_shuffle[6200];
    assign key_original[7142] = key_shuffle[8036];
    assign key_original[7141] = key_shuffle[3693];
    assign key_original[7140] = key_shuffle[6177];
    assign key_original[7139] = key_shuffle[4547];
    assign key_original[7138] = key_shuffle[7061];
    assign key_original[7137] = key_shuffle[134];
    assign key_original[7136] = key_shuffle[188];
    assign key_original[7135] = key_shuffle[6370];
    assign key_original[7134] = key_shuffle[5892];
    assign key_original[7133] = key_shuffle[2815];
    assign key_original[7132] = key_shuffle[5028];
    assign key_original[7131] = key_shuffle[6815];
    assign key_original[7130] = key_shuffle[3029];
    assign key_original[7129] = key_shuffle[3203];
    assign key_original[7128] = key_shuffle[2533];
    assign key_original[7127] = key_shuffle[4577];
    assign key_original[7126] = key_shuffle[946];
    assign key_original[7125] = key_shuffle[5556];
    assign key_original[7124] = key_shuffle[2222];
    assign key_original[7123] = key_shuffle[40];
    assign key_original[7122] = key_shuffle[6375];
    assign key_original[7121] = key_shuffle[5602];
    assign key_original[7120] = key_shuffle[3726];
    assign key_original[7119] = key_shuffle[4881];
    assign key_original[7118] = key_shuffle[1582];
    assign key_original[7117] = key_shuffle[324];
    assign key_original[7116] = key_shuffle[6639];
    assign key_original[7115] = key_shuffle[3389];
    assign key_original[7114] = key_shuffle[5290];
    assign key_original[7113] = key_shuffle[483];
    assign key_original[7112] = key_shuffle[7256];
    assign key_original[7111] = key_shuffle[708];
    assign key_original[7110] = key_shuffle[7551];
    assign key_original[7109] = key_shuffle[5769];
    assign key_original[7108] = key_shuffle[5473];
    assign key_original[7107] = key_shuffle[6612];
    assign key_original[7106] = key_shuffle[616];
    assign key_original[7105] = key_shuffle[8100];
    assign key_original[7104] = key_shuffle[6728];
    assign key_original[7103] = key_shuffle[5988];
    assign key_original[7102] = key_shuffle[2896];
    assign key_original[7101] = key_shuffle[316];
    assign key_original[7100] = key_shuffle[3122];
    assign key_original[7099] = key_shuffle[5325];
    assign key_original[7098] = key_shuffle[1747];
    assign key_original[7097] = key_shuffle[7485];
    assign key_original[7096] = key_shuffle[1320];
    assign key_original[7095] = key_shuffle[1376];
    assign key_original[7094] = key_shuffle[2416];
    assign key_original[7093] = key_shuffle[8179];
    assign key_original[7092] = key_shuffle[7540];
    assign key_original[7091] = key_shuffle[8104];
    assign key_original[7090] = key_shuffle[5090];
    assign key_original[7089] = key_shuffle[4062];
    assign key_original[7088] = key_shuffle[1284];
    assign key_original[7087] = key_shuffle[5469];
    assign key_original[7086] = key_shuffle[5818];
    assign key_original[7085] = key_shuffle[5789];
    assign key_original[7084] = key_shuffle[2870];
    assign key_original[7083] = key_shuffle[2185];
    assign key_original[7082] = key_shuffle[7667];
    assign key_original[7081] = key_shuffle[547];
    assign key_original[7080] = key_shuffle[310];
    assign key_original[7079] = key_shuffle[3606];
    assign key_original[7078] = key_shuffle[1632];
    assign key_original[7077] = key_shuffle[2554];
    assign key_original[7076] = key_shuffle[7231];
    assign key_original[7075] = key_shuffle[5809];
    assign key_original[7074] = key_shuffle[6191];
    assign key_original[7073] = key_shuffle[3087];
    assign key_original[7072] = key_shuffle[352];
    assign key_original[7071] = key_shuffle[5141];
    assign key_original[7070] = key_shuffle[2426];
    assign key_original[7069] = key_shuffle[3];
    assign key_original[7068] = key_shuffle[2872];
    assign key_original[7067] = key_shuffle[6367];
    assign key_original[7066] = key_shuffle[4502];
    assign key_original[7065] = key_shuffle[875];
    assign key_original[7064] = key_shuffle[5518];
    assign key_original[7063] = key_shuffle[4641];
    assign key_original[7062] = key_shuffle[2375];
    assign key_original[7061] = key_shuffle[7763];
    assign key_original[7060] = key_shuffle[6746];
    assign key_original[7059] = key_shuffle[4612];
    assign key_original[7058] = key_shuffle[3955];
    assign key_original[7057] = key_shuffle[1842];
    assign key_original[7056] = key_shuffle[5383];
    assign key_original[7055] = key_shuffle[1542];
    assign key_original[7054] = key_shuffle[1855];
    assign key_original[7053] = key_shuffle[1779];
    assign key_original[7052] = key_shuffle[5743];
    assign key_original[7051] = key_shuffle[678];
    assign key_original[7050] = key_shuffle[1959];
    assign key_original[7049] = key_shuffle[4053];
    assign key_original[7048] = key_shuffle[3563];
    assign key_original[7047] = key_shuffle[4171];
    assign key_original[7046] = key_shuffle[3724];
    assign key_original[7045] = key_shuffle[3082];
    assign key_original[7044] = key_shuffle[5832];
    assign key_original[7043] = key_shuffle[5126];
    assign key_original[7042] = key_shuffle[2801];
    assign key_original[7041] = key_shuffle[6811];
    assign key_original[7040] = key_shuffle[6905];
    assign key_original[7039] = key_shuffle[3034];
    assign key_original[7038] = key_shuffle[6158];
    assign key_original[7037] = key_shuffle[7328];
    assign key_original[7036] = key_shuffle[907];
    assign key_original[7035] = key_shuffle[3893];
    assign key_original[7034] = key_shuffle[6089];
    assign key_original[7033] = key_shuffle[5];
    assign key_original[7032] = key_shuffle[201];
    assign key_original[7031] = key_shuffle[6809];
    assign key_original[7030] = key_shuffle[7117];
    assign key_original[7029] = key_shuffle[7472];
    assign key_original[7028] = key_shuffle[514];
    assign key_original[7027] = key_shuffle[4509];
    assign key_original[7026] = key_shuffle[7894];
    assign key_original[7025] = key_shuffle[1750];
    assign key_original[7024] = key_shuffle[3268];
    assign key_original[7023] = key_shuffle[5084];
    assign key_original[7022] = key_shuffle[6959];
    assign key_original[7021] = key_shuffle[4927];
    assign key_original[7020] = key_shuffle[1269];
    assign key_original[7019] = key_shuffle[5828];
    assign key_original[7018] = key_shuffle[5183];
    assign key_original[7017] = key_shuffle[5036];
    assign key_original[7016] = key_shuffle[3701];
    assign key_original[7015] = key_shuffle[1510];
    assign key_original[7014] = key_shuffle[3491];
    assign key_original[7013] = key_shuffle[853];
    assign key_original[7012] = key_shuffle[6257];
    assign key_original[7011] = key_shuffle[3008];
    assign key_original[7010] = key_shuffle[8161];
    assign key_original[7009] = key_shuffle[2757];
    assign key_original[7008] = key_shuffle[3078];
    assign key_original[7007] = key_shuffle[1914];
    assign key_original[7006] = key_shuffle[1484];
    assign key_original[7005] = key_shuffle[2108];
    assign key_original[7004] = key_shuffle[7360];
    assign key_original[7003] = key_shuffle[3017];
    assign key_original[7002] = key_shuffle[7832];
    assign key_original[7001] = key_shuffle[2702];
    assign key_original[7000] = key_shuffle[102];
    assign key_original[6999] = key_shuffle[465];
    assign key_original[6998] = key_shuffle[2076];
    assign key_original[6997] = key_shuffle[576];
    assign key_original[6996] = key_shuffle[2659];
    assign key_original[6995] = key_shuffle[6836];
    assign key_original[6994] = key_shuffle[1734];
    assign key_original[6993] = key_shuffle[6197];
    assign key_original[6992] = key_shuffle[1834];
    assign key_original[6991] = key_shuffle[5107];
    assign key_original[6990] = key_shuffle[6901];
    assign key_original[6989] = key_shuffle[4580];
    assign key_original[6988] = key_shuffle[125];
    assign key_original[6987] = key_shuffle[6944];
    assign key_original[6986] = key_shuffle[1199];
    assign key_original[6985] = key_shuffle[2445];
    assign key_original[6984] = key_shuffle[5622];
    assign key_original[6983] = key_shuffle[2762];
    assign key_original[6982] = key_shuffle[1073];
    assign key_original[6981] = key_shuffle[5069];
    assign key_original[6980] = key_shuffle[7777];
    assign key_original[6979] = key_shuffle[3702];
    assign key_original[6978] = key_shuffle[5616];
    assign key_original[6977] = key_shuffle[2433];
    assign key_original[6976] = key_shuffle[1975];
    assign key_original[6975] = key_shuffle[4411];
    assign key_original[6974] = key_shuffle[1545];
    assign key_original[6973] = key_shuffle[772];
    assign key_original[6972] = key_shuffle[4403];
    assign key_original[6971] = key_shuffle[4181];
    assign key_original[6970] = key_shuffle[6927];
    assign key_original[6969] = key_shuffle[7727];
    assign key_original[6968] = key_shuffle[1622];
    assign key_original[6967] = key_shuffle[5959];
    assign key_original[6966] = key_shuffle[7891];
    assign key_original[6965] = key_shuffle[3850];
    assign key_original[6964] = key_shuffle[5856];
    assign key_original[6963] = key_shuffle[6428];
    assign key_original[6962] = key_shuffle[4554];
    assign key_original[6961] = key_shuffle[5199];
    assign key_original[6960] = key_shuffle[3367];
    assign key_original[6959] = key_shuffle[4205];
    assign key_original[6958] = key_shuffle[5986];
    assign key_original[6957] = key_shuffle[1678];
    assign key_original[6956] = key_shuffle[6661];
    assign key_original[6955] = key_shuffle[4207];
    assign key_original[6954] = key_shuffle[6328];
    assign key_original[6953] = key_shuffle[6114];
    assign key_original[6952] = key_shuffle[1];
    assign key_original[6951] = key_shuffle[1802];
    assign key_original[6950] = key_shuffle[3490];
    assign key_original[6949] = key_shuffle[18];
    assign key_original[6948] = key_shuffle[1731];
    assign key_original[6947] = key_shuffle[3422];
    assign key_original[6946] = key_shuffle[3009];
    assign key_original[6945] = key_shuffle[6761];
    assign key_original[6944] = key_shuffle[8025];
    assign key_original[6943] = key_shuffle[6917];
    assign key_original[6942] = key_shuffle[4897];
    assign key_original[6941] = key_shuffle[1771];
    assign key_original[6940] = key_shuffle[179];
    assign key_original[6939] = key_shuffle[922];
    assign key_original[6938] = key_shuffle[1393];
    assign key_original[6937] = key_shuffle[7690];
    assign key_original[6936] = key_shuffle[1562];
    assign key_original[6935] = key_shuffle[2615];
    assign key_original[6934] = key_shuffle[140];
    assign key_original[6933] = key_shuffle[6634];
    assign key_original[6932] = key_shuffle[4833];
    assign key_original[6931] = key_shuffle[4839];
    assign key_original[6930] = key_shuffle[4980];
    assign key_original[6929] = key_shuffle[3427];
    assign key_original[6928] = key_shuffle[7114];
    assign key_original[6927] = key_shuffle[3204];
    assign key_original[6926] = key_shuffle[122];
    assign key_original[6925] = key_shuffle[4396];
    assign key_original[6924] = key_shuffle[207];
    assign key_original[6923] = key_shuffle[3909];
    assign key_original[6922] = key_shuffle[3738];
    assign key_original[6921] = key_shuffle[5086];
    assign key_original[6920] = key_shuffle[1999];
    assign key_original[6919] = key_shuffle[7825];
    assign key_original[6918] = key_shuffle[7097];
    assign key_original[6917] = key_shuffle[4477];
    assign key_original[6916] = key_shuffle[4343];
    assign key_original[6915] = key_shuffle[3696];
    assign key_original[6914] = key_shuffle[3011];
    assign key_original[6913] = key_shuffle[1396];
    assign key_original[6912] = key_shuffle[2248];
    assign key_original[6911] = key_shuffle[5801];
    assign key_original[6910] = key_shuffle[7614];
    assign key_original[6909] = key_shuffle[1163];
    assign key_original[6908] = key_shuffle[7636];
    assign key_original[6907] = key_shuffle[4856];
    assign key_original[6906] = key_shuffle[1141];
    assign key_original[6905] = key_shuffle[6221];
    assign key_original[6904] = key_shuffle[3280];
    assign key_original[6903] = key_shuffle[4717];
    assign key_original[6902] = key_shuffle[3995];
    assign key_original[6901] = key_shuffle[2228];
    assign key_original[6900] = key_shuffle[471];
    assign key_original[6899] = key_shuffle[1148];
    assign key_original[6898] = key_shuffle[197];
    assign key_original[6897] = key_shuffle[4327];
    assign key_original[6896] = key_shuffle[3711];
    assign key_original[6895] = key_shuffle[7455];
    assign key_original[6894] = key_shuffle[1843];
    assign key_original[6893] = key_shuffle[1867];
    assign key_original[6892] = key_shuffle[5582];
    assign key_original[6891] = key_shuffle[1997];
    assign key_original[6890] = key_shuffle[6573];
    assign key_original[6889] = key_shuffle[4114];
    assign key_original[6888] = key_shuffle[1744];
    assign key_original[6887] = key_shuffle[3002];
    assign key_original[6886] = key_shuffle[7197];
    assign key_original[6885] = key_shuffle[604];
    assign key_original[6884] = key_shuffle[1317];
    assign key_original[6883] = key_shuffle[3613];
    assign key_original[6882] = key_shuffle[5933];
    assign key_original[6881] = key_shuffle[2994];
    assign key_original[6880] = key_shuffle[746];
    assign key_original[6879] = key_shuffle[5357];
    assign key_original[6878] = key_shuffle[4364];
    assign key_original[6877] = key_shuffle[5054];
    assign key_original[6876] = key_shuffle[7694];
    assign key_original[6875] = key_shuffle[7957];
    assign key_original[6874] = key_shuffle[21];
    assign key_original[6873] = key_shuffle[3095];
    assign key_original[6872] = key_shuffle[2939];
    assign key_original[6871] = key_shuffle[3162];
    assign key_original[6870] = key_shuffle[459];
    assign key_original[6869] = key_shuffle[7399];
    assign key_original[6868] = key_shuffle[4922];
    assign key_original[6867] = key_shuffle[2831];
    assign key_original[6866] = key_shuffle[7559];
    assign key_original[6865] = key_shuffle[7029];
    assign key_original[6864] = key_shuffle[5122];
    assign key_original[6863] = key_shuffle[6421];
    assign key_original[6862] = key_shuffle[614];
    assign key_original[6861] = key_shuffle[312];
    assign key_original[6860] = key_shuffle[718];
    assign key_original[6859] = key_shuffle[5891];
    assign key_original[6858] = key_shuffle[7425];
    assign key_original[6857] = key_shuffle[5216];
    assign key_original[6856] = key_shuffle[7706];
    assign key_original[6855] = key_shuffle[1683];
    assign key_original[6854] = key_shuffle[7630];
    assign key_original[6853] = key_shuffle[3579];
    assign key_original[6852] = key_shuffle[7516];
    assign key_original[6851] = key_shuffle[3765];
    assign key_original[6850] = key_shuffle[5558];
    assign key_original[6849] = key_shuffle[7435];
    assign key_original[6848] = key_shuffle[1349];
    assign key_original[6847] = key_shuffle[3290];
    assign key_original[6846] = key_shuffle[2061];
    assign key_original[6845] = key_shuffle[5146];
    assign key_original[6844] = key_shuffle[6804];
    assign key_original[6843] = key_shuffle[4009];
    assign key_original[6842] = key_shuffle[291];
    assign key_original[6841] = key_shuffle[2696];
    assign key_original[6840] = key_shuffle[3670];
    assign key_original[6839] = key_shuffle[6157];
    assign key_original[6838] = key_shuffle[1818];
    assign key_original[6837] = key_shuffle[7113];
    assign key_original[6836] = key_shuffle[4289];
    assign key_original[6835] = key_shuffle[6239];
    assign key_original[6834] = key_shuffle[1058];
    assign key_original[6833] = key_shuffle[7581];
    assign key_original[6832] = key_shuffle[3891];
    assign key_original[6831] = key_shuffle[1144];
    assign key_original[6830] = key_shuffle[874];
    assign key_original[6829] = key_shuffle[4507];
    assign key_original[6828] = key_shuffle[4064];
    assign key_original[6827] = key_shuffle[755];
    assign key_original[6826] = key_shuffle[3510];
    assign key_original[6825] = key_shuffle[3345];
    assign key_original[6824] = key_shuffle[7009];
    assign key_original[6823] = key_shuffle[4155];
    assign key_original[6822] = key_shuffle[2213];
    assign key_original[6821] = key_shuffle[4112];
    assign key_original[6820] = key_shuffle[6826];
    assign key_original[6819] = key_shuffle[5438];
    assign key_original[6818] = key_shuffle[1701];
    assign key_original[6817] = key_shuffle[2168];
    assign key_original[6816] = key_shuffle[2992];
    assign key_original[6815] = key_shuffle[2578];
    assign key_original[6814] = key_shuffle[566];
    assign key_original[6813] = key_shuffle[4648];
    assign key_original[6812] = key_shuffle[6098];
    assign key_original[6811] = key_shuffle[6730];
    assign key_original[6810] = key_shuffle[7537];
    assign key_original[6809] = key_shuffle[3125];
    assign key_original[6808] = key_shuffle[3450];
    assign key_original[6807] = key_shuffle[7010];
    assign key_original[6806] = key_shuffle[2552];
    assign key_original[6805] = key_shuffle[6117];
    assign key_original[6804] = key_shuffle[6193];
    assign key_original[6803] = key_shuffle[2078];
    assign key_original[6802] = key_shuffle[4383];
    assign key_original[6801] = key_shuffle[2595];
    assign key_original[6800] = key_shuffle[3144];
    assign key_original[6799] = key_shuffle[7089];
    assign key_original[6798] = key_shuffle[4244];
    assign key_original[6797] = key_shuffle[7842];
    assign key_original[6796] = key_shuffle[625];
    assign key_original[6795] = key_shuffle[3771];
    assign key_original[6794] = key_shuffle[7679];
    assign key_original[6793] = key_shuffle[3015];
    assign key_original[6792] = key_shuffle[4262];
    assign key_original[6791] = key_shuffle[290];
    assign key_original[6790] = key_shuffle[3036];
    assign key_original[6789] = key_shuffle[7159];
    assign key_original[6788] = key_shuffle[2680];
    assign key_original[6787] = key_shuffle[1195];
    assign key_original[6786] = key_shuffle[1335];
    assign key_original[6785] = key_shuffle[2195];
    assign key_original[6784] = key_shuffle[5349];
    assign key_original[6783] = key_shuffle[2704];
    assign key_original[6782] = key_shuffle[5760];
    assign key_original[6781] = key_shuffle[6643];
    assign key_original[6780] = key_shuffle[1748];
    assign key_original[6779] = key_shuffle[359];
    assign key_original[6778] = key_shuffle[2996];
    assign key_original[6777] = key_shuffle[6525];
    assign key_original[6776] = key_shuffle[2333];
    assign key_original[6775] = key_shuffle[6829];
    assign key_original[6774] = key_shuffle[5754];
    assign key_original[6773] = key_shuffle[5834];
    assign key_original[6772] = key_shuffle[4965];
    assign key_original[6771] = key_shuffle[2944];
    assign key_original[6770] = key_shuffle[4261];
    assign key_original[6769] = key_shuffle[2904];
    assign key_original[6768] = key_shuffle[2504];
    assign key_original[6767] = key_shuffle[3719];
    assign key_original[6766] = key_shuffle[2354];
    assign key_original[6765] = key_shuffle[4734];
    assign key_original[6764] = key_shuffle[7890];
    assign key_original[6763] = key_shuffle[7535];
    assign key_original[6762] = key_shuffle[6863];
    assign key_original[6761] = key_shuffle[2306];
    assign key_original[6760] = key_shuffle[3472];
    assign key_original[6759] = key_shuffle[1344];
    assign key_original[6758] = key_shuffle[1817];
    assign key_original[6757] = key_shuffle[6878];
    assign key_original[6756] = key_shuffle[1052];
    assign key_original[6755] = key_shuffle[7520];
    assign key_original[6754] = key_shuffle[1374];
    assign key_original[6753] = key_shuffle[8029];
    assign key_original[6752] = key_shuffle[5851];
    assign key_original[6751] = key_shuffle[7753];
    assign key_original[6750] = key_shuffle[6339];
    assign key_original[6749] = key_shuffle[6511];
    assign key_original[6748] = key_shuffle[373];
    assign key_original[6747] = key_shuffle[2331];
    assign key_original[6746] = key_shuffle[1753];
    assign key_original[6745] = key_shuffle[6877];
    assign key_original[6744] = key_shuffle[5796];
    assign key_original[6743] = key_shuffle[1043];
    assign key_original[6742] = key_shuffle[4313];
    assign key_original[6741] = key_shuffle[2644];
    assign key_original[6740] = key_shuffle[89];
    assign key_original[6739] = key_shuffle[227];
    assign key_original[6738] = key_shuffle[2454];
    assign key_original[6737] = key_shuffle[2523];
    assign key_original[6736] = key_shuffle[1807];
    assign key_original[6735] = key_shuffle[2320];
    assign key_original[6734] = key_shuffle[5829];
    assign key_original[6733] = key_shuffle[2952];
    assign key_original[6732] = key_shuffle[1574];
    assign key_original[6731] = key_shuffle[1784];
    assign key_original[6730] = key_shuffle[6052];
    assign key_original[6729] = key_shuffle[6493];
    assign key_original[6728] = key_shuffle[1488];
    assign key_original[6727] = key_shuffle[2843];
    assign key_original[6726] = key_shuffle[8111];
    assign key_original[6725] = key_shuffle[3267];
    assign key_original[6724] = key_shuffle[486];
    assign key_original[6723] = key_shuffle[8068];
    assign key_original[6722] = key_shuffle[3991];
    assign key_original[6721] = key_shuffle[5001];
    assign key_original[6720] = key_shuffle[3302];
    assign key_original[6719] = key_shuffle[5245];
    assign key_original[6718] = key_shuffle[4203];
    assign key_original[6717] = key_shuffle[997];
    assign key_original[6716] = key_shuffle[2875];
    assign key_original[6715] = key_shuffle[92];
    assign key_original[6714] = key_shuffle[2897];
    assign key_original[6713] = key_shuffle[6440];
    assign key_original[6712] = key_shuffle[7652];
    assign key_original[6711] = key_shuffle[1066];
    assign key_original[6710] = key_shuffle[3342];
    assign key_original[6709] = key_shuffle[6475];
    assign key_original[6708] = key_shuffle[4995];
    assign key_original[6707] = key_shuffle[2139];
    assign key_original[6706] = key_shuffle[5385];
    assign key_original[6705] = key_shuffle[4143];
    assign key_original[6704] = key_shuffle[3773];
    assign key_original[6703] = key_shuffle[5472];
    assign key_original[6702] = key_shuffle[5687];
    assign key_original[6701] = key_shuffle[2550];
    assign key_original[6700] = key_shuffle[3173];
    assign key_original[6699] = key_shuffle[6272];
    assign key_original[6698] = key_shuffle[5215];
    assign key_original[6697] = key_shuffle[4533];
    assign key_original[6696] = key_shuffle[6699];
    assign key_original[6695] = key_shuffle[6682];
    assign key_original[6694] = key_shuffle[5857];
    assign key_original[6693] = key_shuffle[1850];
    assign key_original[6692] = key_shuffle[3304];
    assign key_original[6691] = key_shuffle[399];
    assign key_original[6690] = key_shuffle[1427];
    assign key_original[6689] = key_shuffle[610];
    assign key_original[6688] = key_shuffle[2453];
    assign key_original[6687] = key_shuffle[3497];
    assign key_original[6686] = key_shuffle[2058];
    assign key_original[6685] = key_shuffle[7491];
    assign key_original[6684] = key_shuffle[52];
    assign key_original[6683] = key_shuffle[3762];
    assign key_original[6682] = key_shuffle[6388];
    assign key_original[6681] = key_shuffle[462];
    assign key_original[6680] = key_shuffle[401];
    assign key_original[6679] = key_shuffle[2438];
    assign key_original[6678] = key_shuffle[6094];
    assign key_original[6677] = key_shuffle[4830];
    assign key_original[6676] = key_shuffle[132];
    assign key_original[6675] = key_shuffle[852];
    assign key_original[6674] = key_shuffle[4685];
    assign key_original[6673] = key_shuffle[5348];
    assign key_original[6672] = key_shuffle[4491];
    assign key_original[6671] = key_shuffle[1617];
    assign key_original[6670] = key_shuffle[6947];
    assign key_original[6669] = key_shuffle[196];
    assign key_original[6668] = key_shuffle[3752];
    assign key_original[6667] = key_shuffle[10];
    assign key_original[6666] = key_shuffle[5591];
    assign key_original[6665] = key_shuffle[2883];
    assign key_original[6664] = key_shuffle[3619];
    assign key_original[6663] = key_shuffle[6182];
    assign key_original[6662] = key_shuffle[382];
    assign key_original[6661] = key_shuffle[1256];
    assign key_original[6660] = key_shuffle[7741];
    assign key_original[6659] = key_shuffle[3735];
    assign key_original[6658] = key_shuffle[5475];
    assign key_original[6657] = key_shuffle[5994];
    assign key_original[6656] = key_shuffle[7859];
    assign key_original[6655] = key_shuffle[5190];
    assign key_original[6654] = key_shuffle[168];
    assign key_original[6653] = key_shuffle[1476];
    assign key_original[6652] = key_shuffle[6923];
    assign key_original[6651] = key_shuffle[464];
    assign key_original[6650] = key_shuffle[2528];
    assign key_original[6649] = key_shuffle[5077];
    assign key_original[6648] = key_shuffle[7628];
    assign key_original[6647] = key_shuffle[2698];
    assign key_original[6646] = key_shuffle[720];
    assign key_original[6645] = key_shuffle[8075];
    assign key_original[6644] = key_shuffle[5831];
    assign key_original[6643] = key_shuffle[7998];
    assign key_original[6642] = key_shuffle[2301];
    assign key_original[6641] = key_shuffle[2945];
    assign key_original[6640] = key_shuffle[5316];
    assign key_original[6639] = key_shuffle[6081];
    assign key_original[6638] = key_shuffle[7995];
    assign key_original[6637] = key_shuffle[2633];
    assign key_original[6636] = key_shuffle[782];
    assign key_original[6635] = key_shuffle[7503];
    assign key_original[6634] = key_shuffle[3090];
    assign key_original[6633] = key_shuffle[3922];
    assign key_original[6632] = key_shuffle[3842];
    assign key_original[6631] = key_shuffle[1566];
    assign key_original[6630] = key_shuffle[2969];
    assign key_original[6629] = key_shuffle[1904];
    assign key_original[6628] = key_shuffle[4873];
    assign key_original[6627] = key_shuffle[6389];
    assign key_original[6626] = key_shuffle[2837];
    assign key_original[6625] = key_shuffle[2854];
    assign key_original[6624] = key_shuffle[6734];
    assign key_original[6623] = key_shuffle[5545];
    assign key_original[6622] = key_shuffle[3245];
    assign key_original[6621] = key_shuffle[4377];
    assign key_original[6620] = key_shuffle[2964];
    assign key_original[6619] = key_shuffle[482];
    assign key_original[6618] = key_shuffle[4872];
    assign key_original[6617] = key_shuffle[1218];
    assign key_original[6616] = key_shuffle[2075];
    assign key_original[6615] = key_shuffle[3632];
    assign key_original[6614] = key_shuffle[1400];
    assign key_original[6613] = key_shuffle[2795];
    assign key_original[6612] = key_shuffle[328];
    assign key_original[6611] = key_shuffle[7116];
    assign key_original[6610] = key_shuffle[5350];
    assign key_original[6609] = key_shuffle[4500];
    assign key_original[6608] = key_shuffle[3751];
    assign key_original[6607] = key_shuffle[3524];
    assign key_original[6606] = key_shuffle[6817];
    assign key_original[6605] = key_shuffle[7158];
    assign key_original[6604] = key_shuffle[6301];
    assign key_original[6603] = key_shuffle[3733];
    assign key_original[6602] = key_shuffle[3102];
    assign key_original[6601] = key_shuffle[203];
    assign key_original[6600] = key_shuffle[5815];
    assign key_original[6599] = key_shuffle[1935];
    assign key_original[6598] = key_shuffle[4134];
    assign key_original[6597] = key_shuffle[4851];
    assign key_original[6596] = key_shuffle[5617];
    assign key_original[6595] = key_shuffle[5256];
    assign key_original[6594] = key_shuffle[5496];
    assign key_original[6593] = key_shuffle[3281];
    assign key_original[6592] = key_shuffle[2622];
    assign key_original[6591] = key_shuffle[5811];
    assign key_original[6590] = key_shuffle[5970];
    assign key_original[6589] = key_shuffle[6707];
    assign key_original[6588] = key_shuffle[1980];
    assign key_original[6587] = key_shuffle[3688];
    assign key_original[6586] = key_shuffle[524];
    assign key_original[6585] = key_shuffle[6973];
    assign key_original[6584] = key_shuffle[7768];
    assign key_original[6583] = key_shuffle[1880];
    assign key_original[6582] = key_shuffle[1482];
    assign key_original[6581] = key_shuffle[6966];
    assign key_original[6580] = key_shuffle[2967];
    assign key_original[6579] = key_shuffle[5521];
    assign key_original[6578] = key_shuffle[4326];
    assign key_original[6577] = key_shuffle[1183];
    assign key_original[6576] = key_shuffle[4276];
    assign key_original[6575] = key_shuffle[632];
    assign key_original[6574] = key_shuffle[7647];
    assign key_original[6573] = key_shuffle[4871];
    assign key_original[6572] = key_shuffle[3152];
    assign key_original[6571] = key_shuffle[6977];
    assign key_original[6570] = key_shuffle[6663];
    assign key_original[6569] = key_shuffle[2321];
    assign key_original[6568] = key_shuffle[5601];
    assign key_original[6567] = key_shuffle[1724];
    assign key_original[6566] = key_shuffle[7400];
    assign key_original[6565] = key_shuffle[58];
    assign key_original[6564] = key_shuffle[7127];
    assign key_original[6563] = key_shuffle[6860];
    assign key_original[6562] = key_shuffle[5498];
    assign key_original[6561] = key_shuffle[5702];
    assign key_original[6560] = key_shuffle[4721];
    assign key_original[6559] = key_shuffle[1700];
    assign key_original[6558] = key_shuffle[692];
    assign key_original[6557] = key_shuffle[3448];
    assign key_original[6556] = key_shuffle[7078];
    assign key_original[6555] = key_shuffle[618];
    assign key_original[6554] = key_shuffle[5441];
    assign key_original[6553] = key_shuffle[3038];
    assign key_original[6552] = key_shuffle[4816];
    assign key_original[6551] = key_shuffle[42];
    assign key_original[6550] = key_shuffle[8058];
    assign key_original[6549] = key_shuffle[914];
    assign key_original[6548] = key_shuffle[1089];
    assign key_original[6547] = key_shuffle[2727];
    assign key_original[6546] = key_shuffle[893];
    assign key_original[6545] = key_shuffle[3094];
    assign key_original[6544] = key_shuffle[7];
    assign key_original[6543] = key_shuffle[6206];
    assign key_original[6542] = key_shuffle[6551];
    assign key_original[6541] = key_shuffle[5719];
    assign key_original[6540] = key_shuffle[6925];
    assign key_original[6539] = key_shuffle[176];
    assign key_original[6538] = key_shuffle[5427];
    assign key_original[6537] = key_shuffle[829];
    assign key_original[6536] = key_shuffle[2556];
    assign key_original[6535] = key_shuffle[913];
    assign key_original[6534] = key_shuffle[538];
    assign key_original[6533] = key_shuffle[2292];
    assign key_original[6532] = key_shuffle[3411];
    assign key_original[6531] = key_shuffle[980];
    assign key_original[6530] = key_shuffle[1598];
    assign key_original[6529] = key_shuffle[8144];
    assign key_original[6528] = key_shuffle[5944];
    assign key_original[6527] = key_shuffle[3967];
    assign key_original[6526] = key_shuffle[8082];
    assign key_original[6525] = key_shuffle[4158];
    assign key_original[6524] = key_shuffle[5233];
    assign key_original[6523] = key_shuffle[2082];
    assign key_original[6522] = key_shuffle[2155];
    assign key_original[6521] = key_shuffle[1286];
    assign key_original[6520] = key_shuffle[1267];
    assign key_original[6519] = key_shuffle[5224];
    assign key_original[6518] = key_shuffle[6801];
    assign key_original[6517] = key_shuffle[6608];
    assign key_original[6516] = key_shuffle[7469];
    assign key_original[6515] = key_shuffle[3347];
    assign key_original[6514] = key_shuffle[2197];
    assign key_original[6513] = key_shuffle[7111];
    assign key_original[6512] = key_shuffle[4079];
    assign key_original[6511] = key_shuffle[6592];
    assign key_original[6510] = key_shuffle[6943];
    assign key_original[6509] = key_shuffle[2613];
    assign key_original[6508] = key_shuffle[4880];
    assign key_original[6507] = key_shuffle[5361];
    assign key_original[6506] = key_shuffle[1714];
    assign key_original[6505] = key_shuffle[728];
    assign key_original[6504] = key_shuffle[7571];
    assign key_original[6503] = key_shuffle[3539];
    assign key_original[6502] = key_shuffle[2389];
    assign key_original[6501] = key_shuffle[208];
    assign key_original[6500] = key_shuffle[157];
    assign key_original[6499] = key_shuffle[2474];
    assign key_original[6498] = key_shuffle[4536];
    assign key_original[6497] = key_shuffle[6251];
    assign key_original[6496] = key_shuffle[6467];
    assign key_original[6495] = key_shuffle[1514];
    assign key_original[6494] = key_shuffle[4492];
    assign key_original[6493] = key_shuffle[2866];
    assign key_original[6492] = key_shuffle[8102];
    assign key_original[6491] = key_shuffle[2879];
    assign key_original[6490] = key_shuffle[1227];
    assign key_original[6489] = key_shuffle[519];
    assign key_original[6488] = key_shuffle[2806];
    assign key_original[6487] = key_shuffle[4296];
    assign key_original[6486] = key_shuffle[2890];
    assign key_original[6485] = key_shuffle[5305];
    assign key_original[6484] = key_shuffle[2586];
    assign key_original[6483] = key_shuffle[2350];
    assign key_original[6482] = key_shuffle[7077];
    assign key_original[6481] = key_shuffle[2716];
    assign key_original[6480] = key_shuffle[4608];
    assign key_original[6479] = key_shuffle[6599];
    assign key_original[6478] = key_shuffle[4041];
    assign key_original[6477] = key_shuffle[5289];
    assign key_original[6476] = key_shuffle[3254];
    assign key_original[6475] = key_shuffle[1262];
    assign key_original[6474] = key_shuffle[4543];
    assign key_original[6473] = key_shuffle[2824];
    assign key_original[6472] = key_shuffle[2707];
    assign key_original[6471] = key_shuffle[756];
    assign key_original[6470] = key_shuffle[4138];
    assign key_original[6469] = key_shuffle[6530];
    assign key_original[6468] = key_shuffle[7674];
    assign key_original[6467] = key_shuffle[1246];
    assign key_original[6466] = key_shuffle[6381];
    assign key_original[6465] = key_shuffle[3879];
    assign key_original[6464] = key_shuffle[2326];
    assign key_original[6463] = key_shuffle[1675];
    assign key_original[6462] = key_shuffle[3359];
    assign key_original[6461] = key_shuffle[5159];
    assign key_original[6460] = key_shuffle[2774];
    assign key_original[6459] = key_shuffle[3885];
    assign key_original[6458] = key_shuffle[2720];
    assign key_original[6457] = key_shuffle[7885];
    assign key_original[6456] = key_shuffle[7668];
    assign key_original[6455] = key_shuffle[8013];
    assign key_original[6454] = key_shuffle[4441];
    assign key_original[6453] = key_shuffle[2961];
    assign key_original[6452] = key_shuffle[5530];
    assign key_original[6451] = key_shuffle[7532];
    assign key_original[6450] = key_shuffle[2792];
    assign key_original[6449] = key_shuffle[4986];
    assign key_original[6448] = key_shuffle[7437];
    assign key_original[6447] = key_shuffle[1070];
    assign key_original[6446] = key_shuffle[7880];
    assign key_original[6445] = key_shuffle[4286];
    assign key_original[6444] = key_shuffle[5189];
    assign key_original[6443] = key_shuffle[80];
    assign key_original[6442] = key_shuffle[972];
    assign key_original[6441] = key_shuffle[6235];
    assign key_original[6440] = key_shuffle[1800];
    assign key_original[6439] = key_shuffle[2599];
    assign key_original[6438] = key_shuffle[702];
    assign key_original[6437] = key_shuffle[421];
    assign key_original[6436] = key_shuffle[3823];
    assign key_original[6435] = key_shuffle[7931];
    assign key_original[6434] = key_shuffle[7306];
    assign key_original[6433] = key_shuffle[3760];
    assign key_original[6432] = key_shuffle[6396];
    assign key_original[6431] = key_shuffle[3037];
    assign key_original[6430] = key_shuffle[1826];
    assign key_original[6429] = key_shuffle[6310];
    assign key_original[6428] = key_shuffle[1856];
    assign key_original[6427] = key_shuffle[6990];
    assign key_original[6426] = key_shuffle[4370];
    assign key_original[6425] = key_shuffle[2421];
    assign key_original[6424] = key_shuffle[2052];
    assign key_original[6423] = key_shuffle[6791];
    assign key_original[6422] = key_shuffle[1629];
    assign key_original[6421] = key_shuffle[4243];
    assign key_original[6420] = key_shuffle[724];
    assign key_original[6419] = key_shuffle[3511];
    assign key_original[6418] = key_shuffle[2793];
    assign key_original[6417] = key_shuffle[3467];
    assign key_original[6416] = key_shuffle[527];
    assign key_original[6415] = key_shuffle[7059];
    assign key_original[6414] = key_shuffle[1181];
    assign key_original[6413] = key_shuffle[4273];
    assign key_original[6412] = key_shuffle[8146];
    assign key_original[6411] = key_shuffle[640];
    assign key_original[6410] = key_shuffle[8170];
    assign key_original[6409] = key_shuffle[882];
    assign key_original[6408] = key_shuffle[5896];
    assign key_original[6407] = key_shuffle[4918];
    assign key_original[6406] = key_shuffle[273];
    assign key_original[6405] = key_shuffle[3261];
    assign key_original[6404] = key_shuffle[6092];
    assign key_original[6403] = key_shuffle[911];
    assign key_original[6402] = key_shuffle[7883];
    assign key_original[6401] = key_shuffle[791];
    assign key_original[6400] = key_shuffle[3882];
    assign key_original[6399] = key_shuffle[578];
    assign key_original[6398] = key_shuffle[6725];
    assign key_original[6397] = key_shuffle[2404];
    assign key_original[6396] = key_shuffle[5494];
    assign key_original[6395] = key_shuffle[7253];
    assign key_original[6394] = key_shuffle[5858];
    assign key_original[6393] = key_shuffle[4843];
    assign key_original[6392] = key_shuffle[4541];
    assign key_original[6391] = key_shuffle[5382];
    assign key_original[6390] = key_shuffle[6470];
    assign key_original[6389] = key_shuffle[4065];
    assign key_original[6388] = key_shuffle[3133];
    assign key_original[6387] = key_shuffle[700];
    assign key_original[6386] = key_shuffle[1011];
    assign key_original[6385] = key_shuffle[2811];
    assign key_original[6384] = key_shuffle[6224];
    assign key_original[6383] = key_shuffle[5938];
    assign key_original[6382] = key_shuffle[1830];
    assign key_original[6381] = key_shuffle[6557];
    assign key_original[6380] = key_shuffle[4926];
    assign key_original[6379] = key_shuffle[2186];
    assign key_original[6378] = key_shuffle[2848];
    assign key_original[6377] = key_shuffle[6026];
    assign key_original[6376] = key_shuffle[215];
    assign key_original[6375] = key_shuffle[2498];
    assign key_original[6374] = key_shuffle[5952];
    assign key_original[6373] = key_shuffle[1243];
    assign key_original[6372] = key_shuffle[4671];
    assign key_original[6371] = key_shuffle[7866];
    assign key_original[6370] = key_shuffle[7238];
    assign key_original[6369] = key_shuffle[5669];
    assign key_original[6368] = key_shuffle[2216];
    assign key_original[6367] = key_shuffle[1124];
    assign key_original[6366] = key_shuffle[7168];
    assign key_original[6365] = key_shuffle[7489];
    assign key_original[6364] = key_shuffle[3307];
    assign key_original[6363] = key_shuffle[7284];
    assign key_original[6362] = key_shuffle[6986];
    assign key_original[6361] = key_shuffle[3700];
    assign key_original[6360] = key_shuffle[4760];
    assign key_original[6359] = key_shuffle[3927];
    assign key_original[6358] = key_shuffle[8017];
    assign key_original[6357] = key_shuffle[596];
    assign key_original[6356] = key_shuffle[6140];
    assign key_original[6355] = key_shuffle[5087];
    assign key_original[6354] = key_shuffle[1272];
    assign key_original[6353] = key_shuffle[5660];
    assign key_original[6352] = key_shuffle[374];
    assign key_original[6351] = key_shuffle[1039];
    assign key_original[6350] = key_shuffle[7884];
    assign key_original[6349] = key_shuffle[2397];
    assign key_original[6348] = key_shuffle[4805];
    assign key_original[6347] = key_shuffle[6134];
    assign key_original[6346] = key_shuffle[3534];
    assign key_original[6345] = key_shuffle[371];
    assign key_original[6344] = key_shuffle[3118];
    assign key_original[6343] = key_shuffle[3071];
    assign key_original[6342] = key_shuffle[3778];
    assign key_original[6341] = key_shuffle[5276];
    assign key_original[6340] = key_shuffle[516];
    assign key_original[6339] = key_shuffle[6178];
    assign key_original[6338] = key_shuffle[2895];
    assign key_original[6337] = key_shuffle[7258];
    assign key_original[6336] = key_shuffle[552];
    assign key_original[6335] = key_shuffle[2274];
    assign key_original[6334] = key_shuffle[288];
    assign key_original[6333] = key_shuffle[199];
    assign key_original[6332] = key_shuffle[5730];
    assign key_original[6331] = key_shuffle[246];
    assign key_original[6330] = key_shuffle[7038];
    assign key_original[6329] = key_shuffle[2304];
    assign key_original[6328] = key_shuffle[5943];
    assign key_original[6327] = key_shuffle[6362];
    assign key_original[6326] = key_shuffle[2286];
    assign key_original[6325] = key_shuffle[3802];
    assign key_original[6324] = key_shuffle[7709];
    assign key_original[6323] = key_shuffle[487];
    assign key_original[6322] = key_shuffle[4495];
    assign key_original[6321] = key_shuffle[7564];
    assign key_original[6320] = key_shuffle[3241];
    assign key_original[6319] = key_shuffle[1528];
    assign key_original[6318] = key_shuffle[6244];
    assign key_original[6317] = key_shuffle[6124];
    assign key_original[6316] = key_shuffle[8];
    assign key_original[6315] = key_shuffle[7391];
    assign key_original[6314] = key_shuffle[3820];
    assign key_original[6313] = key_shuffle[225];
    assign key_original[6312] = key_shuffle[8041];
    assign key_original[6311] = key_shuffle[508];
    assign key_original[6310] = key_shuffle[6874];
    assign key_original[6309] = key_shuffle[3535];
    assign key_original[6308] = key_shuffle[5654];
    assign key_original[6307] = key_shuffle[1537];
    assign key_original[6306] = key_shuffle[24];
    assign key_original[6305] = key_shuffle[2518];
    assign key_original[6304] = key_shuffle[5042];
    assign key_original[6303] = key_shuffle[726];
    assign key_original[6302] = key_shuffle[1864];
    assign key_original[6301] = key_shuffle[4444];
    assign key_original[6300] = key_shuffle[5600];
    assign key_original[6299] = key_shuffle[410];
    assign key_original[6298] = key_shuffle[1074];
    assign key_original[6297] = key_shuffle[7632];
    assign key_original[6296] = key_shuffle[6088];
    assign key_original[6295] = key_shuffle[2791];
    assign key_original[6294] = key_shuffle[6903];
    assign key_original[6293] = key_shuffle[6930];
    assign key_original[6292] = key_shuffle[5318];
    assign key_original[6291] = key_shuffle[7230];
    assign key_original[6290] = key_shuffle[4545];
    assign key_original[6289] = key_shuffle[8076];
    assign key_original[6288] = key_shuffle[2860];
    assign key_original[6287] = key_shuffle[2759];
    assign key_original[6286] = key_shuffle[6093];
    assign key_original[6285] = key_shuffle[3523];
    assign key_original[6284] = key_shuffle[683];
    assign key_original[6283] = key_shuffle[198];
    assign key_original[6282] = key_shuffle[194];
    assign key_original[6281] = key_shuffle[5063];
    assign key_original[6280] = key_shuffle[3656];
    assign key_original[6279] = key_shuffle[2923];
    assign key_original[6278] = key_shuffle[4683];
    assign key_original[6277] = key_shuffle[1394];
    assign key_original[6276] = key_shuffle[7362];
    assign key_original[6275] = key_shuffle[6256];
    assign key_original[6274] = key_shuffle[6722];
    assign key_original[6273] = key_shuffle[1912];
    assign key_original[6272] = key_shuffle[7137];
    assign key_original[6271] = key_shuffle[2849];
    assign key_original[6270] = key_shuffle[456];
    assign key_original[6269] = key_shuffle[3966];
    assign key_original[6268] = key_shuffle[2583];
    assign key_original[6267] = key_shuffle[3083];
    assign key_original[6266] = key_shuffle[5534];
    assign key_original[6265] = key_shuffle[5898];
    assign key_original[6264] = key_shuffle[3236];
    assign key_original[6263] = key_shuffle[6786];
    assign key_original[6262] = key_shuffle[6347];
    assign key_original[6261] = key_shuffle[4693];
    assign key_original[6260] = key_shuffle[1590];
    assign key_original[6259] = key_shuffle[387];
    assign key_original[6258] = key_shuffle[338];
    assign key_original[6257] = key_shuffle[2668];
    assign key_original[6256] = key_shuffle[3665];
    assign key_original[6255] = key_shuffle[1251];
    assign key_original[6254] = key_shuffle[1548];
    assign key_original[6253] = key_shuffle[5167];
    assign key_original[6252] = key_shuffle[2918];
    assign key_original[6251] = key_shuffle[2347];
    assign key_original[6250] = key_shuffle[1938];
    assign key_original[6249] = key_shuffle[8185];
    assign key_original[6248] = key_shuffle[1947];
    assign key_original[6247] = key_shuffle[3892];
    assign key_original[6246] = key_shuffle[5022];
    assign key_original[6245] = key_shuffle[2544];
    assign key_original[6244] = key_shuffle[8101];
    assign key_original[6243] = key_shuffle[3496];
    assign key_original[6242] = key_shuffle[6409];
    assign key_original[6241] = key_shuffle[896];
    assign key_original[6240] = key_shuffle[3033];
    assign key_original[6239] = key_shuffle[7641];
    assign key_original[6238] = key_shuffle[792];
    assign key_original[6237] = key_shuffle[4757];
    assign key_original[6236] = key_shuffle[6776];
    assign key_original[6235] = key_shuffle[3950];
    assign key_original[6234] = key_shuffle[2934];
    assign key_original[6233] = key_shuffle[1763];
    assign key_original[6232] = key_shuffle[7700];
    assign key_original[6231] = key_shuffle[6297];
    assign key_original[6230] = key_shuffle[706];
    assign key_original[6229] = key_shuffle[7319];
    assign key_original[6228] = key_shuffle[6866];
    assign key_original[6227] = key_shuffle[3513];
    assign key_original[6226] = key_shuffle[4714];
    assign key_original[6225] = key_shuffle[3158];
    assign key_original[6224] = key_shuffle[5508];
    assign key_original[6223] = key_shuffle[5726];
    assign key_original[6222] = key_shuffle[3843];
    assign key_original[6221] = key_shuffle[1160];
    assign key_original[6220] = key_shuffle[4800];
    assign key_original[6219] = key_shuffle[3767];
    assign key_original[6218] = key_shuffle[4097];
    assign key_original[6217] = key_shuffle[1336];
    assign key_original[6216] = key_shuffle[318];
    assign key_original[6215] = key_shuffle[7899];
    assign key_original[6214] = key_shuffle[7326];
    assign key_original[6213] = key_shuffle[4682];
    assign key_original[6212] = key_shuffle[6993];
    assign key_original[6211] = key_shuffle[3540];
    assign key_original[6210] = key_shuffle[732];
    assign key_original[6209] = key_shuffle[5571];
    assign key_original[6208] = key_shuffle[5552];
    assign key_original[6207] = key_shuffle[1984];
    assign key_original[6206] = key_shuffle[6788];
    assign key_original[6205] = key_shuffle[2368];
    assign key_original[6204] = key_shuffle[8081];
    assign key_original[6203] = key_shuffle[7785];
    assign key_original[6202] = key_shuffle[773];
    assign key_original[6201] = key_shuffle[7509];
    assign key_original[6200] = key_shuffle[697];
    assign key_original[6199] = key_shuffle[5279];
    assign key_original[6198] = key_shuffle[4164];
    assign key_original[6197] = key_shuffle[7611];
    assign key_original[6196] = key_shuffle[6430];
    assign key_original[6195] = key_shuffle[1235];
    assign key_original[6194] = key_shuffle[819];
    assign key_original[6193] = key_shuffle[5745];
    assign key_original[6192] = key_shuffle[7067];
    assign key_original[6191] = key_shuffle[5578];
    assign key_original[6190] = key_shuffle[3819];
    assign key_original[6189] = key_shuffle[5166];
    assign key_original[6188] = key_shuffle[6284];
    assign key_original[6187] = key_shuffle[4110];
    assign key_original[6186] = key_shuffle[7858];
    assign key_original[6185] = key_shuffle[6220];
    assign key_original[6184] = key_shuffle[1131];
    assign key_original[6183] = key_shuffle[3140];
    assign key_original[6182] = key_shuffle[7441];
    assign key_original[6181] = key_shuffle[6056];
    assign key_original[6180] = key_shuffle[5206];
    assign key_original[6179] = key_shuffle[130];
    assign key_original[6178] = key_shuffle[3500];
    assign key_original[6177] = key_shuffle[584];
    assign key_original[6176] = key_shuffle[1464];
    assign key_original[6175] = key_shuffle[7347];
    assign key_original[6174] = key_shuffle[4841];
    assign key_original[6173] = key_shuffle[531];
    assign key_original[6172] = key_shuffle[4912];
    assign key_original[6171] = key_shuffle[65];
    assign key_original[6170] = key_shuffle[6647];
    assign key_original[6169] = key_shuffle[1757];
    assign key_original[6168] = key_shuffle[1328];
    assign key_original[6167] = key_shuffle[4340];
    assign key_original[6166] = key_shuffle[4768];
    assign key_original[6165] = key_shuffle[2745];
    assign key_original[6164] = key_shuffle[4499];
    assign key_original[6163] = key_shuffle[536];
    assign key_original[6162] = key_shuffle[780];
    assign key_original[6161] = key_shuffle[1170];
    assign key_original[6160] = key_shuffle[64];
    assign key_original[6159] = key_shuffle[7203];
    assign key_original[6158] = key_shuffle[6890];
    assign key_original[6157] = key_shuffle[4005];
    assign key_original[6156] = key_shuffle[869];
    assign key_original[6155] = key_shuffle[3785];
    assign key_original[6154] = key_shuffle[4855];
    assign key_original[6153] = key_shuffle[7954];
    assign key_original[6152] = key_shuffle[6108];
    assign key_original[6151] = key_shuffle[7255];
    assign key_original[6150] = key_shuffle[7024];
    assign key_original[6149] = key_shuffle[2662];
    assign key_original[6148] = key_shuffle[3603];
    assign key_original[6147] = key_shuffle[3180];
    assign key_original[6146] = key_shuffle[5513];
    assign key_original[6145] = key_shuffle[2294];
    assign key_original[6144] = key_shuffle[1847];
    assign key_original[6143] = key_shuffle[4515];
    assign key_original[6142] = key_shuffle[790];
    assign key_original[6141] = key_shuffle[7940];
    assign key_original[6140] = key_shuffle[4689];
    assign key_original[6139] = key_shuffle[3106];
    assign key_original[6138] = key_shuffle[7278];
    assign key_original[6137] = key_shuffle[4631];
    assign key_original[6136] = key_shuffle[2047];
    assign key_original[6135] = key_shuffle[4393];
    assign key_original[6134] = key_shuffle[1083];
    assign key_original[6133] = key_shuffle[6752];
    assign key_original[6132] = key_shuffle[6775];
    assign key_original[6131] = key_shuffle[5467];
    assign key_original[6130] = key_shuffle[804];
    assign key_original[6129] = key_shuffle[6512];
    assign key_original[6128] = key_shuffle[5049];
    assign key_original[6127] = key_shuffle[7394];
    assign key_original[6126] = key_shuffle[7914];
    assign key_original[6125] = key_shuffle[1721];
    assign key_original[6124] = key_shuffle[3310];
    assign key_original[6123] = key_shuffle[173];
    assign key_original[6122] = key_shuffle[3589];
    assign key_original[6121] = key_shuffle[2154];
    assign key_original[6120] = key_shuffle[3402];
    assign key_original[6119] = key_shuffle[7561];
    assign key_original[6118] = key_shuffle[2677];
    assign key_original[6117] = key_shuffle[4222];
    assign key_original[6116] = key_shuffle[4801];
    assign key_original[6115] = key_shuffle[5538];
    assign key_original[6114] = key_shuffle[4644];
    assign key_original[6113] = key_shuffle[6165];
    assign key_original[6112] = key_shuffle[830];
    assign key_original[6111] = key_shuffle[332];
    assign key_original[6110] = key_shuffle[6883];
    assign key_original[6109] = key_shuffle[5737];
    assign key_original[6108] = key_shuffle[474];
    assign key_original[6107] = key_shuffle[79];
    assign key_original[6106] = key_shuffle[3551];
    assign key_original[6105] = key_shuffle[2589];
    assign key_original[6104] = key_shuffle[3908];
    assign key_original[6103] = key_shuffle[1892];
    assign key_original[6102] = key_shuffle[3697];
    assign key_original[6101] = key_shuffle[3270];
    assign key_original[6100] = key_shuffle[3601];
    assign key_original[6099] = key_shuffle[5132];
    assign key_original[6098] = key_shuffle[4542];
    assign key_original[6097] = key_shuffle[4910];
    assign key_original[6096] = key_shuffle[1242];
    assign key_original[6095] = key_shuffle[4350];
    assign key_original[6094] = key_shuffle[2280];
    assign key_original[6093] = key_shuffle[4621];
    assign key_original[6092] = key_shuffle[2775];
    assign key_original[6091] = key_shuffle[7456];
    assign key_original[6090] = key_shuffle[7961];
    assign key_original[6089] = key_shuffle[3965];
    assign key_original[6088] = key_shuffle[2183];
    assign key_original[6087] = key_shuffle[654];
    assign key_original[6086] = key_shuffle[1241];
    assign key_original[6085] = key_shuffle[2768];
    assign key_original[6084] = key_shuffle[837];
    assign key_original[6083] = key_shuffle[3024];
    assign key_original[6082] = key_shuffle[4960];
    assign key_original[6081] = key_shuffle[3883];
    assign key_original[6080] = key_shuffle[2114];
    assign key_original[6079] = key_shuffle[4268];
    assign key_original[6078] = key_shuffle[5095];
    assign key_original[6077] = key_shuffle[6099];
    assign key_original[6076] = key_shuffle[2681];
    assign key_original[6075] = key_shuffle[2434];
    assign key_original[6074] = key_shuffle[5968];
    assign key_original[6073] = key_shuffle[2922];
    assign key_original[6072] = key_shuffle[4100];
    assign key_original[6071] = key_shuffle[636];
    assign key_original[6070] = key_shuffle[1258];
    assign key_original[6069] = key_shuffle[6252];
    assign key_original[6068] = key_shuffle[4359];
    assign key_original[6067] = key_shuffle[4788];
    assign key_original[6066] = key_shuffle[5064];
    assign key_original[6065] = key_shuffle[2217];
    assign key_original[6064] = key_shuffle[7375];
    assign key_original[6063] = key_shuffle[5100];
    assign key_original[6062] = key_shuffle[5218];
    assign key_original[6061] = key_shuffle[4940];
    assign key_original[6060] = key_shuffle[5824];
    assign key_original[6059] = key_shuffle[988];
    assign key_original[6058] = key_shuffle[1762];
    assign key_original[6057] = key_shuffle[5002];
    assign key_original[6056] = key_shuffle[3275];
    assign key_original[6055] = key_shuffle[3754];
    assign key_original[6054] = key_shuffle[5684];
    assign key_original[6053] = key_shuffle[6255];
    assign key_original[6052] = key_shuffle[2505];
    assign key_original[6051] = key_shuffle[6552];
    assign key_original[6050] = key_shuffle[2738];
    assign key_original[6049] = key_shuffle[7098];
    assign key_original[6048] = key_shuffle[3732];
    assign key_original[6047] = key_shuffle[2122];
    assign key_original[6046] = key_shuffle[6824];
    assign key_original[6045] = key_shuffle[5260];
    assign key_original[6044] = key_shuffle[7244];
    assign key_original[6043] = key_shuffle[7605];
    assign key_original[6042] = key_shuffle[6001];
    assign key_original[6041] = key_shuffle[649];
    assign key_original[6040] = key_shuffle[1307];
    assign key_original[6039] = key_shuffle[442];
    assign key_original[6038] = key_shuffle[7022];
    assign key_original[6037] = key_shuffle[7464];
    assign key_original[6036] = key_shuffle[1226];
    assign key_original[6035] = key_shuffle[7019];
    assign key_original[6034] = key_shuffle[3982];
    assign key_original[6033] = key_shuffle[3946];
    assign key_original[6032] = key_shuffle[3548];
    assign key_original[6031] = key_shuffle[7069];
    assign key_original[6030] = key_shuffle[1560];
    assign key_original[6029] = key_shuffle[6377];
    assign key_original[6028] = key_shuffle[2314];
    assign key_original[6027] = key_shuffle[4250];
    assign key_original[6026] = key_shuffle[1413];
    assign key_original[6025] = key_shuffle[1592];
    assign key_original[6024] = key_shuffle[1061];
    assign key_original[6023] = key_shuffle[2661];
    assign key_original[6022] = key_shuffle[5517];
    assign key_original[6021] = key_shuffle[5025];
    assign key_original[6020] = key_shuffle[6309];
    assign key_original[6019] = key_shuffle[4699];
    assign key_original[6018] = key_shuffle[3640];
    assign key_original[6017] = key_shuffle[3265];
    assign key_original[6016] = key_shuffle[7035];
    assign key_original[6015] = key_shuffle[2508];
    assign key_original[6014] = key_shuffle[5605];
    assign key_original[6013] = key_shuffle[6142];
    assign key_original[6012] = key_shuffle[428];
    assign key_original[6011] = key_shuffle[2987];
    assign key_original[6010] = key_shuffle[3353];
    assign key_original[6009] = key_shuffle[2778];
    assign key_original[6008] = key_shuffle[3303];
    assign key_original[6007] = key_shuffle[5982];
    assign key_original[6006] = key_shuffle[119];
    assign key_original[6005] = key_shuffle[0];
    assign key_original[6004] = key_shuffle[7817];
    assign key_original[6003] = key_shuffle[5148];
    assign key_original[6002] = key_shuffle[1475];
    assign key_original[6001] = key_shuffle[7750];
    assign key_original[6000] = key_shuffle[4342];
    assign key_original[5999] = key_shuffle[2431];
    assign key_original[5998] = key_shuffle[3315];
    assign key_original[5997] = key_shuffle[193];
    assign key_original[5996] = key_shuffle[7703];
    assign key_original[5995] = key_shuffle[1795];
    assign key_original[5994] = key_shuffle[6072];
    assign key_original[5993] = key_shuffle[7685];
    assign key_original[5992] = key_shuffle[3705];
    assign key_original[5991] = key_shuffle[165];
    assign key_original[5990] = key_shuffle[6680];
    assign key_original[5989] = key_shuffle[920];
    assign key_original[5988] = key_shuffle[441];
    assign key_original[5987] = key_shuffle[394];
    assign key_original[5986] = key_shuffle[4845];
    assign key_original[5985] = key_shuffle[1502];
    assign key_original[5984] = key_shuffle[4552];
    assign key_original[5983] = key_shuffle[6213];
    assign key_original[5982] = key_shuffle[1416];
    assign key_original[5981] = key_shuffle[5875];
    assign key_original[5980] = key_shuffle[1007];
    assign key_original[5979] = key_shuffle[1786];
    assign key_original[5978] = key_shuffle[4704];
    assign key_original[5977] = key_shuffle[1766];
    assign key_original[5976] = key_shuffle[7810];
    assign key_original[5975] = key_shuffle[2959];
    assign key_original[5974] = key_shuffle[7000];
    assign key_original[5973] = key_shuffle[2832];
    assign key_original[5972] = key_shuffle[2128];
    assign key_original[5971] = key_shuffle[7594];
    assign key_original[5970] = key_shuffle[5990];
    assign key_original[5969] = key_shuffle[1943];
    assign key_original[5968] = key_shuffle[3676];
    assign key_original[5967] = key_shuffle[5093];
    assign key_original[5966] = key_shuffle[6303];
    assign key_original[5965] = key_shuffle[7847];
    assign key_original[5964] = key_shuffle[1024];
    assign key_original[5963] = key_shuffle[303];
    assign key_original[5962] = key_shuffle[7980];
    assign key_original[5961] = key_shuffle[7656];
    assign key_original[5960] = key_shuffle[2300];
    assign key_original[5959] = key_shuffle[6032];
    assign key_original[5958] = key_shuffle[4373];
    assign key_original[5957] = key_shuffle[4847];
    assign key_original[5956] = key_shuffle[3098];
    assign key_original[5955] = key_shuffle[7927];
    assign key_original[5954] = key_shuffle[4388];
    assign key_original[5953] = key_shuffle[6956];
    assign key_original[5952] = key_shuffle[2231];
    assign key_original[5951] = key_shuffle[7192];
    assign key_original[5950] = key_shuffle[989];
    assign key_original[5949] = key_shuffle[4535];
    assign key_original[5948] = key_shuffle[7575];
    assign key_original[5947] = key_shuffle[269];
    assign key_original[5946] = key_shuffle[4645];
    assign key_original[5945] = key_shuffle[4642];
    assign key_original[5944] = key_shuffle[7812];
    assign key_original[5943] = key_shuffle[4368];
    assign key_original[5942] = key_shuffle[3063];
    assign key_original[5941] = key_shuffle[7661];
    assign key_original[5940] = key_shuffle[1648];
    assign key_original[5939] = key_shuffle[3866];
    assign key_original[5938] = key_shuffle[3372];
    assign key_original[5937] = key_shuffle[94];
    assign key_original[5936] = key_shuffle[5926];
    assign key_original[5935] = key_shuffle[8110];
    assign key_original[5934] = key_shuffle[4522];
    assign key_original[5933] = key_shuffle[1038];
    assign key_original[5932] = key_shuffle[292];
    assign key_original[5931] = key_shuffle[7984];
    assign key_original[5930] = key_shuffle[8014];
    assign key_original[5929] = key_shuffle[6263];
    assign key_original[5928] = key_shuffle[3723];
    assign key_original[5927] = key_shuffle[6657];
    assign key_original[5926] = key_shuffle[7148];
    assign key_original[5925] = key_shuffle[1085];
    assign key_original[5924] = key_shuffle[2448];
    assign key_original[5923] = key_shuffle[3923];
    assign key_original[5922] = key_shuffle[4779];
    assign key_original[5921] = key_shuffle[1467];
    assign key_original[5920] = key_shuffle[2223];
    assign key_original[5919] = key_shuffle[5031];
    assign key_original[5918] = key_shuffle[5400];
    assign key_original[5917] = key_shuffle[1260];
    assign key_original[5916] = key_shuffle[7839];
    assign key_original[5915] = key_shuffle[5454];
    assign key_original[5914] = key_shuffle[5979];
    assign key_original[5913] = key_shuffle[1945];
    assign key_original[5912] = key_shuffle[7865];
    assign key_original[5911] = key_shuffle[6483];
    assign key_original[5910] = key_shuffle[3393];
    assign key_original[5909] = key_shuffle[5599];
    assign key_original[5908] = key_shuffle[3833];
    assign key_original[5907] = key_shuffle[305];
    assign key_original[5906] = key_shuffle[3952];
    assign key_original[5905] = key_shuffle[936];
    assign key_original[5904] = key_shuffle[5401];
    assign key_original[5903] = key_shuffle[1441];
    assign key_original[5902] = key_shuffle[7963];
    assign key_original[5901] = key_shuffle[867];
    assign key_original[5900] = key_shuffle[429];
    assign key_original[5899] = key_shuffle[6839];
    assign key_original[5898] = key_shuffle[4319];
    assign key_original[5897] = key_shuffle[3568];
    assign key_original[5896] = key_shuffle[6410];
    assign key_original[5895] = key_shuffle[2830];
    assign key_original[5894] = key_shuffle[7265];
    assign key_original[5893] = key_shuffle[6210];
    assign key_original[5892] = key_shuffle[3777];
    assign key_original[5891] = key_shuffle[3206];
    assign key_original[5890] = key_shuffle[5932];
    assign key_original[5889] = key_shuffle[2995];
    assign key_original[5888] = key_shuffle[849];
    assign key_original[5887] = key_shuffle[8044];
    assign key_original[5886] = key_shuffle[2152];
    assign key_original[5885] = key_shuffle[3248];
    assign key_original[5884] = key_shuffle[7650];
    assign key_original[5883] = key_shuffle[4749];
    assign key_original[5882] = key_shuffle[509];
    assign key_original[5881] = key_shuffle[415];
    assign key_original[5880] = key_shuffle[7841];
    assign key_original[5879] = key_shuffle[546];
    assign key_original[5878] = key_shuffle[7214];
    assign key_original[5877] = key_shuffle[3478];
    assign key_original[5876] = key_shuffle[885];
    assign key_original[5875] = key_shuffle[5615];
    assign key_original[5874] = key_shuffle[3564];
    assign key_original[5873] = key_shuffle[4111];
    assign key_original[5872] = key_shuffle[4540];
    assign key_original[5871] = key_shuffle[6386];
    assign key_original[5870] = key_shuffle[1956];
    assign key_original[5869] = key_shuffle[166];
    assign key_original[5868] = key_shuffle[3997];
    assign key_original[5867] = key_shuffle[4168];
    assign key_original[5866] = key_shuffle[5570];
    assign key_original[5865] = key_shuffle[581];
    assign key_original[5864] = key_shuffle[131];
    assign key_original[5863] = key_shuffle[4513];
    assign key_original[5862] = key_shuffle[3333];
    assign key_original[5861] = key_shuffle[8045];
    assign key_original[5860] = key_shuffle[3430];
    assign key_original[5859] = key_shuffle[5627];
    assign key_original[5858] = key_shuffle[6718];
    assign key_original[5857] = key_shuffle[148];
    assign key_original[5856] = key_shuffle[2588];
    assign key_original[5855] = key_shuffle[4221];
    assign key_original[5854] = key_shuffle[261];
    assign key_original[5853] = key_shuffle[6369];
    assign key_original[5852] = key_shuffle[2856];
    assign key_original[5851] = key_shuffle[2754];
    assign key_original[5850] = key_shuffle[2840];
    assign key_original[5849] = key_shuffle[4988];
    assign key_original[5848] = key_shuffle[4568];
    assign key_original[5847] = key_shuffle[3558];
    assign key_original[5846] = key_shuffle[3799];
    assign key_original[5845] = key_shuffle[2332];
    assign key_original[5844] = key_shuffle[6958];
    assign key_original[5843] = key_shuffle[1071];
    assign key_original[5842] = key_shuffle[8178];
    assign key_original[5841] = key_shuffle[7965];
    assign key_original[5840] = key_shuffle[7478];
    assign key_original[5839] = key_shuffle[4530];
    assign key_original[5838] = key_shuffle[6768];
    assign key_original[5837] = key_shuffle[4553];
    assign key_original[5836] = key_shuffle[3390];
    assign key_original[5835] = key_shuffle[4709];
    assign key_original[5834] = key_shuffle[6779];
    assign key_original[5833] = key_shuffle[3685];
    assign key_original[5832] = key_shuffle[1293];
    assign key_original[5831] = key_shuffle[6975];
    assign key_original[5830] = key_shuffle[2298];
    assign key_original[5829] = key_shuffle[7924];
    assign key_original[5828] = key_shuffle[3003];
    assign key_original[5827] = key_shuffle[4336];
    assign key_original[5826] = key_shuffle[1332];
    assign key_original[5825] = key_shuffle[2512];
    assign key_original[5824] = key_shuffle[5455];
    assign key_original[5823] = key_shuffle[6102];
    assign key_original[5822] = key_shuffle[5776];
    assign key_original[5821] = key_shuffle[6145];
    assign key_original[5820] = key_shuffle[7737];
    assign key_original[5819] = key_shuffle[3928];
    assign key_original[5818] = key_shuffle[383];
    assign key_original[5817] = key_shuffle[6068];
    assign key_original[5816] = key_shuffle[7151];
    assign key_original[5815] = key_shuffle[118];
    assign key_original[5814] = key_shuffle[8083];
    assign key_original[5813] = key_shuffle[2208];
    assign key_original[5812] = key_shuffle[2728];
    assign key_original[5811] = key_shuffle[443];
    assign key_original[5810] = key_shuffle[6954];
    assign key_original[5809] = key_shuffle[973];
    assign key_original[5808] = key_shuffle[3255];
    assign key_original[5807] = key_shuffle[7494];
    assign key_original[5806] = key_shuffle[2119];
    assign key_original[5805] = key_shuffle[6561];
    assign key_original[5804] = key_shuffle[2157];
    assign key_original[5803] = key_shuffle[1259];
    assign key_original[5802] = key_shuffle[3869];
    assign key_original[5801] = key_shuffle[5269];
    assign key_original[5800] = key_shuffle[7738];
    assign key_original[5799] = key_shuffle[4452];
    assign key_original[5798] = key_shuffle[6714];
    assign key_original[5797] = key_shuffle[7637];
    assign key_original[5796] = key_shuffle[7005];
    assign key_original[5795] = key_shuffle[5563];
    assign key_original[5794] = key_shuffle[1576];
    assign key_original[5793] = key_shuffle[7619];
    assign key_original[5792] = key_shuffle[8046];
    assign key_original[5791] = key_shuffle[3545];
    assign key_original[5790] = key_shuffle[2678];
    assign key_original[5789] = key_shuffle[3649];
    assign key_original[5788] = key_shuffle[2261];
    assign key_original[5787] = key_shuffle[6879];
    assign key_original[5786] = key_shuffle[3763];
    assign key_original[5785] = key_shuffle[5655];
    assign key_original[5784] = key_shuffle[1736];
    assign key_original[5783] = key_shuffle[6457];
    assign key_original[5782] = key_shuffle[663];
    assign key_original[5781] = key_shuffle[1463];
    assign key_original[5780] = key_shuffle[7534];
    assign key_original[5779] = key_shuffle[8050];
    assign key_original[5778] = key_shuffle[3791];
    assign key_original[5777] = key_shuffle[7926];
    assign key_original[5776] = key_shuffle[4994];
    assign key_original[5775] = key_shuffle[4321];
    assign key_original[5774] = key_shuffle[4438];
    assign key_original[5773] = key_shuffle[976];
    assign key_original[5772] = key_shuffle[7164];
    assign key_original[5771] = key_shuffle[2534];
    assign key_original[5770] = key_shuffle[6955];
    assign key_original[5769] = key_shuffle[4347];
    assign key_original[5768] = key_shuffle[3730];
    assign key_original[5767] = key_shuffle[4339];
    assign key_original[5766] = key_shuffle[8106];
    assign key_original[5765] = key_shuffle[6232];
    assign key_original[5764] = key_shuffle[7888];
    assign key_original[5763] = key_shuffle[872];
    assign key_original[5762] = key_shuffle[5399];
    assign key_original[5761] = key_shuffle[3538];
    assign key_original[5760] = key_shuffle[7642];
    assign key_original[5759] = key_shuffle[4119];
    assign key_original[5758] = key_shuffle[5478];
    assign key_original[5757] = key_shuffle[9];
    assign key_original[5756] = key_shuffle[121];
    assign key_original[5755] = key_shuffle[3237];
    assign key_original[5754] = key_shuffle[4977];
    assign key_original[5753] = key_shuffle[2221];
    assign key_original[5752] = key_shuffle[1992];
    assign key_original[5751] = key_shuffle[6217];
    assign key_original[5750] = key_shuffle[4144];
    assign key_original[5749] = key_shuffle[5555];
    assign key_original[5748] = key_shuffle[1849];
    assign key_original[5747] = key_shuffle[2073];
    assign key_original[5746] = key_shuffle[729];
    assign key_original[5745] = key_shuffle[2348];
    assign key_original[5744] = key_shuffle[7588];
    assign key_original[5743] = key_shuffle[680];
    assign key_original[5742] = key_shuffle[4068];
    assign key_original[5741] = key_shuffle[31];
    assign key_original[5740] = key_shuffle[5307];
    assign key_original[5739] = key_shuffle[1920];
    assign key_original[5738] = key_shuffle[4941];
    assign key_original[5737] = key_shuffle[626];
    assign key_original[5736] = key_shuffle[924];
    assign key_original[5735] = key_shuffle[6653];
    assign key_original[5734] = key_shuffle[5045];
    assign key_original[5733] = key_shuffle[2499];
    assign key_original[5732] = key_shuffle[6556];
    assign key_original[5731] = key_shuffle[5873];
    assign key_original[5730] = key_shuffle[1030];
    assign key_original[5729] = key_shuffle[6420];
    assign key_original[5728] = key_shuffle[2900];
    assign key_original[5727] = key_shuffle[5452];
    assign key_original[5726] = key_shuffle[6152];
    assign key_original[5725] = key_shuffle[6055];
    assign key_original[5724] = key_shuffle[3864];
    assign key_original[5723] = key_shuffle[2766];
    assign key_original[5722] = key_shuffle[7733];
    assign key_original[5721] = key_shuffle[8074];
    assign key_original[5720] = key_shuffle[1792];
    assign key_original[5719] = key_shuffle[5321];
    assign key_original[5718] = key_shuffle[1681];
    assign key_original[5717] = key_shuffle[3627];
    assign key_original[5716] = key_shuffle[6497];
    assign key_original[5715] = key_shuffle[7161];
    assign key_original[5714] = key_shuffle[6004];
    assign key_original[5713] = key_shuffle[2829];
    assign key_original[5712] = key_shuffle[2531];
    assign key_original[5711] = key_shuffle[146];
    assign key_original[5710] = key_shuffle[3561];
    assign key_original[5709] = key_shuffle[5683];
    assign key_original[5708] = key_shuffle[6238];
    assign key_original[5707] = key_shuffle[6563];
    assign key_original[5706] = key_shuffle[3728];
    assign key_original[5705] = key_shuffle[7546];
    assign key_original[5704] = key_shuffle[7988];
    assign key_original[5703] = key_shuffle[4765];
    assign key_original[5702] = key_shuffle[7282];
    assign key_original[5701] = key_shuffle[5887];
    assign key_original[5700] = key_shuffle[1862];
    assign key_original[5699] = key_shuffle[6357];
    assign key_original[5698] = key_shuffle[3065];
    assign key_original[5697] = key_shuffle[2054];
    assign key_original[5696] = key_shuffle[3234];
    assign key_original[5695] = key_shuffle[1596];
    assign key_original[5694] = key_shuffle[5484];
    assign key_original[5693] = key_shuffle[4505];
    assign key_original[5692] = key_shuffle[1927];
    assign key_original[5691] = key_shuffle[4778];
    assign key_original[5690] = key_shuffle[7856];
    assign key_original[5689] = key_shuffle[1405];
    assign key_original[5688] = key_shuffle[4290];
    assign key_original[5687] = key_shuffle[1121];
    assign key_original[5686] = key_shuffle[1232];
    assign key_original[5685] = key_shuffle[3056];
    assign key_original[5684] = key_shuffle[1410];
    assign key_original[5683] = key_shuffle[2382];
    assign key_original[5682] = key_shuffle[3499];
    assign key_original[5681] = key_shuffle[2763];
    assign key_original[5680] = key_shuffle[4802];
    assign key_original[5679] = key_shuffle[115];
    assign key_original[5678] = key_shuffle[3556];
    assign key_original[5677] = key_shuffle[1430];
    assign key_original[5676] = key_shuffle[3218];
    assign key_original[5675] = key_shuffle[1626];
    assign key_original[5674] = key_shuffle[5753];
    assign key_original[5673] = key_shuffle[774];
    assign key_original[5672] = key_shuffle[5536];
    assign key_original[5671] = key_shuffle[8031];
    assign key_original[5670] = key_shuffle[5750];
    assign key_original[5669] = key_shuffle[6992];
    assign key_original[5668] = key_shuffle[5871];
    assign key_original[5667] = key_shuffle[1871];
    assign key_original[5666] = key_shuffle[3623];
    assign key_original[5665] = key_shuffle[6276];
    assign key_original[5664] = key_shuffle[6223];
    assign key_original[5663] = key_shuffle[5038];
    assign key_original[5662] = key_shuffle[3099];
    assign key_original[5661] = key_shuffle[2802];
    assign key_original[5660] = key_shuffle[7047];
    assign key_original[5659] = key_shuffle[5066];
    assign key_original[5658] = key_shuffle[7978];
    assign key_original[5657] = key_shuffle[6233];
    assign key_original[5656] = key_shuffle[3358];
    assign key_original[5655] = key_shuffle[3266];
    assign key_original[5654] = key_shuffle[337];
    assign key_original[5653] = key_shuffle[321];
    assign key_original[5652] = key_shuffle[3277];
    assign key_original[5651] = key_shuffle[86];
    assign key_original[5650] = key_shuffle[1186];
    assign key_original[5649] = key_shuffle[2190];
    assign key_original[5648] = key_shuffle[5927];
    assign key_original[5647] = key_shuffle[6567];
    assign key_original[5646] = key_shuffle[6982];
    assign key_original[5645] = key_shuffle[665];
    assign key_original[5644] = key_shuffle[6459];
    assign key_original[5643] = key_shuffle[1609];
    assign key_original[5642] = key_shuffle[5037];
    assign key_original[5641] = key_shuffle[7149];
    assign key_original[5640] = key_shuffle[2091];
    assign key_original[5639] = key_shuffle[7367];
    assign key_original[5638] = key_shuffle[765];
    assign key_original[5637] = key_shuffle[5716];
    assign key_original[5636] = key_shuffle[5837];
    assign key_original[5635] = key_shuffle[5608];
    assign key_original[5634] = key_shuffle[1305];
    assign key_original[5633] = key_shuffle[707];
    assign key_original[5632] = key_shuffle[4708];
    assign key_original[5631] = key_shuffle[1278];
    assign key_original[5630] = key_shuffle[2835];
    assign key_original[5629] = key_shuffle[2949];
    assign key_original[5628] = key_shuffle[4353];
    assign key_original[5627] = key_shuffle[7597];
    assign key_original[5626] = key_shuffle[5304];
    assign key_original[5625] = key_shuffle[7967];
    assign key_original[5624] = key_shuffle[6558];
    assign key_original[5623] = key_shuffle[1221];
    assign key_original[5622] = key_shuffle[244];
    assign key_original[5621] = key_shuffle[2919];
    assign key_original[5620] = key_shuffle[7401];
    assign key_original[5619] = key_shuffle[479];
    assign key_original[5618] = key_shuffle[71];
    assign key_original[5617] = key_shuffle[5894];
    assign key_original[5616] = key_shuffle[7237];
    assign key_original[5615] = key_shuffle[5954];
    assign key_original[5614] = key_shuffle[3969];
    assign key_original[5613] = key_shuffle[5142];
    assign key_original[5612] = key_shuffle[4953];
    assign key_original[5611] = key_shuffle[2220];
    assign key_original[5610] = key_shuffle[985];
    assign key_original[5609] = key_shuffle[1523];
    assign key_original[5608] = key_shuffle[5326];
    assign key_original[5607] = key_shuffle[3745];
    assign key_original[5606] = key_shuffle[6820];
    assign key_original[5605] = key_shuffle[930];
    assign key_original[5604] = key_shuffle[3257];
    assign key_original[5603] = key_shuffle[2857];
    assign key_original[5602] = key_shuffle[2756];
    assign key_original[5601] = key_shuffle[8079];
    assign key_original[5600] = key_shuffle[339];
    assign key_original[5599] = key_shuffle[1571];
    assign key_original[5598] = key_shuffle[7458];
    assign key_original[5597] = key_shuffle[7786];
    assign key_original[5596] = key_shuffle[1657];
    assign key_original[5595] = key_shuffle[507];
    assign key_original[5594] = key_shuffle[4519];
    assign key_original[5593] = key_shuffle[3546];
    assign key_original[5592] = key_shuffle[4294];
    assign key_original[5591] = key_shuffle[6038];
    assign key_original[5590] = key_shuffle[5434];
    assign key_original[5589] = key_shuffle[917];
    assign key_original[5588] = key_shuffle[7349];
    assign key_original[5587] = key_shuffle[6488];
    assign key_original[5586] = key_shuffle[189];
    assign key_original[5585] = key_shuffle[212];
    assign key_original[5584] = key_shuffle[1162];
    assign key_original[5583] = key_shuffle[661];
    assign key_original[5582] = key_shuffle[634];
    assign key_original[5581] = key_shuffle[4137];
    assign key_original[5580] = key_shuffle[247];
    assign key_original[5579] = key_shuffle[4606];
    assign key_original[5578] = key_shuffle[7048];
    assign key_original[5577] = key_shuffle[1013];
    assign key_original[5576] = key_shuffle[1970];
    assign key_original[5575] = key_shuffle[2640];
    assign key_original[5574] = key_shuffle[7816];
    assign key_original[5573] = key_shuffle[6794];
    assign key_original[5572] = key_shuffle[6192];
    assign key_original[5571] = key_shuffle[5461];
    assign key_original[5570] = key_shuffle[3080];
    assign key_original[5569] = key_shuffle[5656];
    assign key_original[5568] = key_shuffle[8132];
    assign key_original[5567] = key_shuffle[1188];
    assign key_original[5566] = key_shuffle[7639];
    assign key_original[5565] = key_shuffle[6589];
    assign key_original[5564] = key_shuffle[7488];
    assign key_original[5563] = key_shuffle[4822];
    assign key_original[5562] = key_shuffle[1965];
    assign key_original[5561] = key_shuffle[4458];
    assign key_original[5560] = key_shuffle[4651];
    assign key_original[5559] = key_shuffle[2572];
    assign key_original[5558] = key_shuffle[948];
    assign key_original[5557] = key_shuffle[4297];
    assign key_original[5556] = key_shuffle[1767];
    assign key_original[5555] = key_shuffle[7872];
    assign key_original[5554] = key_shuffle[2247];
    assign key_original[5553] = key_shuffle[7951];
    assign key_original[5552] = key_shuffle[5120];
    assign key_original[5551] = key_shuffle[2166];
    assign key_original[5550] = key_shuffle[283];
    assign key_original[5549] = key_shuffle[580];
    assign key_original[5548] = key_shuffle[6553];
    assign key_original[5547] = key_shuffle[7781];
    assign key_original[5546] = key_shuffle[1477];
    assign key_original[5545] = key_shuffle[6859];
    assign key_original[5544] = key_shuffle[8048];
    assign key_original[5543] = key_shuffle[5758];
    assign key_original[5542] = key_shuffle[4748];
    assign key_original[5541] = key_shuffle[7001];
    assign key_original[5540] = key_shuffle[3780];
    assign key_original[5539] = key_shuffle[7294];
    assign key_original[5538] = key_shuffle[4966];
    assign key_original[5537] = key_shuffle[4124];
    assign key_original[5536] = key_shuffle[5236];
    assign key_original[5535] = key_shuffle[7734];
    assign key_original[5534] = key_shuffle[4764];
    assign key_original[5533] = key_shuffle[4389];
    assign key_original[5532] = key_shuffle[529];
    assign key_original[5531] = key_shuffle[903];
    assign key_original[5530] = key_shuffle[2145];
    assign key_original[5529] = key_shuffle[2105];
    assign key_original[5528] = key_shuffle[3250];
    assign key_original[5527] = key_shuffle[565];
    assign key_original[5526] = key_shuffle[1950];
    assign key_original[5525] = key_shuffle[5859];
    assign key_original[5524] = key_shuffle[977];
    assign key_original[5523] = key_shuffle[1285];
    assign key_original[5522] = key_shuffle[6503];
    assign key_original[5521] = key_shuffle[5625];
    assign key_original[5520] = key_shuffle[6230];
    assign key_original[5519] = key_shuffle[3171];
    assign key_original[5518] = key_shuffle[4496];
    assign key_original[5517] = key_shuffle[2638];
    assign key_original[5516] = key_shuffle[6841];
    assign key_original[5515] = key_shuffle[1570];
    assign key_original[5514] = key_shuffle[6679];
    assign key_original[5513] = key_shuffle[6387];
    assign key_original[5512] = key_shuffle[6593];
    assign key_original[5511] = key_shuffle[3041];
    assign key_original[5510] = key_shuffle[4162];
    assign key_original[5509] = key_shuffle[8123];
    assign key_original[5508] = key_shuffle[7202];
    assign key_original[5507] = key_shuffle[4448];
    assign key_original[5506] = key_shuffle[6686];
    assign key_original[5505] = key_shuffle[99];
    assign key_original[5504] = key_shuffle[4378];
    assign key_original[5503] = key_shuffle[2366];
    assign key_original[5502] = key_shuffle[2193];
    assign key_original[5501] = key_shuffle[7756];
    assign key_original[5500] = key_shuffle[2447];
    assign key_original[5499] = key_shuffle[7123];
    assign key_original[5498] = key_shuffle[4027];
    assign key_original[5497] = key_shuffle[4357];
    assign key_original[5496] = key_shuffle[1933];
    assign key_original[5495] = key_shuffle[2660];
    assign key_original[5494] = key_shuffle[7115];
    assign key_original[5493] = key_shuffle[6447];
    assign key_original[5492] = key_shuffle[8152];
    assign key_original[5491] = key_shuffle[4975];
    assign key_original[5490] = key_shuffle[2624];
    assign key_original[5489] = key_shuffle[1318];
    assign key_original[5488] = key_shuffle[513];
    assign key_original[5487] = key_shuffle[7717];
    assign key_original[5486] = key_shuffle[6453];
    assign key_original[5485] = key_shuffle[574];
    assign key_original[5484] = key_shuffle[2845];
    assign key_original[5483] = key_shuffle[2827];
    assign key_original[5482] = key_shuffle[2798];
    assign key_original[5481] = key_shuffle[653];
    assign key_original[5480] = key_shuffle[6010];
    assign key_original[5479] = key_shuffle[1534];
    assign key_original[5478] = key_shuffle[4433];
    assign key_original[5477] = key_shuffle[480];
    assign key_original[5476] = key_shuffle[213];
    assign key_original[5475] = key_shuffle[2112];
    assign key_original[5474] = key_shuffle[2656];
    assign key_original[5473] = key_shuffle[6659];
    assign key_original[5472] = key_shuffle[5062];
    assign key_original[5471] = key_shuffle[6665];
    assign key_original[5470] = key_shuffle[2214];
    assign key_original[5469] = key_shuffle[3831];
    assign key_original[5468] = key_shuffle[1062];
    assign key_original[5467] = key_shuffle[7348];
    assign key_original[5466] = key_shuffle[4188];
    assign key_original[5465] = key_shuffle[7153];
    assign key_original[5464] = key_shuffle[1599];
    assign key_original[5463] = key_shuffle[5713];
    assign key_original[5462] = key_shuffle[5453];
    assign key_original[5461] = key_shuffle[7368];
    assign key_original[5460] = key_shuffle[2497];
    assign key_original[5459] = key_shuffle[2752];
    assign key_original[5458] = key_shuffle[3030];
    assign key_original[5457] = key_shuffle[5284];
    assign key_original[5456] = key_shuffle[4429];
    assign key_original[5455] = key_shuffle[7468];
    assign key_original[5454] = key_shuffle[2329];
    assign key_original[5453] = key_shuffle[3934];
    assign key_original[5452] = key_shuffle[7079];
    assign key_original[5451] = key_shuffle[1177];
    assign key_original[5450] = key_shuffle[4583];
    assign key_original[5449] = key_shuffle[957];
    assign key_original[5448] = key_shuffle[1668];
    assign key_original[5447] = key_shuffle[6967];
    assign key_original[5446] = key_shuffle[5372];
    assign key_original[5445] = key_shuffle[469];
    assign key_original[5444] = key_shuffle[4161];
    assign key_original[5443] = key_shuffle[2008];
    assign key_original[5442] = key_shuffle[6040];
    assign key_original[5441] = key_shuffle[5848];
    assign key_original[5440] = key_shuffle[6688];
    assign key_original[5439] = key_shuffle[2784];
    assign key_original[5438] = key_shuffle[7953];
    assign key_original[5437] = key_shuffle[4270];
    assign key_original[5436] = key_shuffle[3537];
    assign key_original[5435] = key_shuffle[4182];
    assign key_original[5434] = key_shuffle[5285];
    assign key_original[5433] = key_shuffle[4532];
    assign key_original[5432] = key_shuffle[1308];
    assign key_original[5431] = key_shuffle[1636];
    assign key_original[5430] = key_shuffle[499];
    assign key_original[5429] = key_shuffle[7302];
    assign key_original[5428] = key_shuffle[7599];
    assign key_original[5427] = key_shuffle[4237];
    assign key_original[5426] = key_shuffle[5989];
    assign key_original[5425] = key_shuffle[3332];
    assign key_original[5424] = key_shuffle[4236];
    assign key_original[5423] = key_shuffle[1176];
    assign key_original[5422] = key_shuffle[5173];
    assign key_original[5421] = key_shuffle[2235];
    assign key_original[5420] = key_shuffle[7937];
    assign key_original[5419] = key_shuffle[757];
    assign key_original[5418] = key_shuffle[1321];
    assign key_original[5417] = key_shuffle[1618];
    assign key_original[5416] = key_shuffle[742];
    assign key_original[5415] = key_shuffle[7312];
    assign key_original[5414] = key_shuffle[413];
    assign key_original[5413] = key_shuffle[4557];
    assign key_original[5412] = key_shuffle[7224];
    assign key_original[5411] = key_shuffle[4597];
    assign key_original[5410] = key_shuffle[7846];
    assign key_original[5409] = key_shuffle[6022];
    assign key_original[5408] = key_shuffle[1531];
    assign key_original[5407] = key_shuffle[2102];
    assign key_original[5406] = key_shuffle[5354];
    assign key_original[5405] = key_shuffle[6581];
    assign key_original[5404] = key_shuffle[4218];
    assign key_original[5403] = key_shuffle[3271];
    assign key_original[5402] = key_shuffle[8141];
    assign key_original[5401] = key_shuffle[3783];
    assign key_original[5400] = key_shuffle[7934];
    assign key_original[5399] = key_shuffle[3880];
    assign key_original[5398] = key_shuffle[6812];
    assign key_original[5397] = key_shuffle[5688];
    assign key_original[5396] = key_shuffle[3214];
    assign key_original[5395] = key_shuffle[7528];
    assign key_original[5394] = key_shuffle[1197];
    assign key_original[5393] = key_shuffle[5041];
    assign key_original[5392] = key_shuffle[6769];
    assign key_original[5391] = key_shuffle[3348];
    assign key_original[5390] = key_shuffle[7558];
    assign key_original[5389] = key_shuffle[6838];
    assign key_original[5388] = key_shuffle[628];
    assign key_original[5387] = key_shuffle[6242];
    assign key_original[5386] = key_shuffle[2269];
    assign key_original[5385] = key_shuffle[1798];
    assign key_original[5384] = key_shuffle[2262];
    assign key_original[5383] = key_shuffle[2786];
    assign key_original[5382] = key_shuffle[4867];
    assign key_original[5381] = key_shuffle[6566];
    assign key_original[5380] = key_shuffle[2600];
    assign key_original[5379] = key_shuffle[3878];
    assign key_original[5378] = key_shuffle[4835];
    assign key_original[5377] = key_shuffle[3830];
    assign key_original[5376] = key_shuffle[7536];
    assign key_original[5375] = key_shuffle[541];
    assign key_original[5374] = key_shuffle[2991];
    assign key_original[5373] = key_shuffle[1381];
    assign key_original[5372] = key_shuffle[1535];
    assign key_original[5371] = key_shuffle[2010];
    assign key_original[5370] = key_shuffle[2734];
    assign key_original[5369] = key_shuffle[6317];
    assign key_original[5368] = key_shuffle[7543];
    assign key_original[5367] = key_shuffle[4204];
    assign key_original[5366] = key_shuffle[7329];
    assign key_original[5365] = key_shuffle[2143];
    assign key_original[5364] = key_shuffle[961];
    assign key_original[5363] = key_shuffle[1159];
    assign key_original[5362] = key_shuffle[4854];
    assign key_original[5361] = key_shuffle[3392];
    assign key_original[5360] = key_shuffle[4213];
    assign key_original[5359] = key_shuffle[1949];
    assign key_original[5358] = key_shuffle[7511];
    assign key_original[5357] = key_shuffle[2187];
    assign key_original[5356] = key_shuffle[6621];
    assign key_original[5355] = key_shuffle[6454];
    assign key_original[5354] = key_shuffle[7204];
    assign key_original[5353] = key_shuffle[856];
    assign key_original[5352] = key_shuffle[695];
    assign key_original[5351] = key_shuffle[7172];
    assign key_original[5350] = key_shuffle[3741];
    assign key_original[5349] = key_shuffle[8043];
    assign key_original[5348] = key_shuffle[6678];
    assign key_original[5347] = key_shuffle[4284];
    assign key_original[5346] = key_shuffle[2914];
    assign key_original[5345] = key_shuffle[2457];
    assign key_original[5344] = key_shuffle[1270];
    assign key_original[5343] = key_shuffle[1200];
    assign key_original[5342] = key_shuffle[5949];
    assign key_original[5341] = key_shuffle[1065];
    assign key_original[5340] = key_shuffle[8149];
    assign key_original[5339] = key_shuffle[5424];
    assign key_original[5338] = key_shuffle[6962];
    assign key_original[5337] = key_shuffle[6431];
    assign key_original[5336] = key_shuffle[7945];
    assign key_original[5335] = key_shuffle[2560];
    assign key_original[5334] = key_shuffle[7490];
    assign key_original[5333] = key_shuffle[1905];
    assign key_original[5332] = key_shuffle[7772];
    assign key_original[5331] = key_shuffle[7790];
    assign key_original[5330] = key_shuffle[6695];
    assign key_original[5329] = key_shuffle[2353];
    assign key_original[5328] = key_shuffle[4152];
    assign key_original[5327] = key_shuffle[5306];
    assign key_original[5326] = key_shuffle[3658];
    assign key_original[5325] = key_shuffle[3731];
    assign key_original[5324] = key_shuffle[6656];
    assign key_original[5323] = key_shuffle[1875];
    assign key_original[5322] = key_shuffle[7243];
    assign key_original[5321] = key_shuffle[1171];
    assign key_original[5320] = key_shuffle[3182];
    assign key_original[5319] = key_shuffle[3594];
    assign key_original[5318] = key_shuffle[8097];
    assign key_original[5317] = key_shuffle[6641];
    assign key_original[5316] = key_shuffle[2469];
    assign key_original[5315] = key_shuffle[3349];
    assign key_original[5314] = key_shuffle[4067];
    assign key_original[5313] = key_shuffle[1020];
    assign key_original[5312] = key_shuffle[1279];
    assign key_original[5311] = key_shuffle[6724];
    assign key_original[5310] = key_shuffle[7334];
    assign key_original[5309] = key_shuffle[1709];
    assign key_original[5308] = key_shuffle[3440];
    assign key_original[5307] = key_shuffle[7498];
    assign key_original[5306] = key_shuffle[3044];
    assign key_original[5305] = key_shuffle[1765];
    assign key_original[5304] = key_shuffle[2200];
    assign key_original[5303] = key_shuffle[1691];
    assign key_original[5302] = key_shuffle[1090];
    assign key_original[5301] = key_shuffle[3356];
    assign key_original[5300] = key_shuffle[560];
    assign key_original[5299] = key_shuffle[2450];
    assign key_original[5298] = key_shuffle[1139];
    assign key_original[5297] = key_shuffle[6871];
    assign key_original[5296] = key_shuffle[2577];
    assign key_original[5295] = key_shuffle[5701];
    assign key_original[5294] = key_shuffle[2901];
    assign key_original[5293] = key_shuffle[7886];
    assign key_original[5292] = key_shuffle[3424];
    assign key_original[5291] = key_shuffle[2511];
    assign key_original[5290] = key_shuffle[1092];
    assign key_original[5289] = key_shuffle[3235];
    assign key_original[5288] = key_shuffle[6189];
    assign key_original[5287] = key_shuffle[7217];
    assign key_original[5286] = key_shuffle[5955];
    assign key_original[5285] = key_shuffle[2403];
    assign key_original[5284] = key_shuffle[1541];
    assign key_original[5283] = key_shuffle[3520];
    assign key_original[5282] = key_shuffle[2169];
    assign key_original[5281] = key_shuffle[3164];
    assign key_original[5280] = key_shuffle[6418];
    assign key_original[5279] = key_shuffle[5791];
    assign key_original[5278] = key_shuffle[4430];
    assign key_original[5277] = key_shuffle[397];
    assign key_original[5276] = key_shuffle[6888];
    assign key_original[5275] = key_shuffle[6462];
    assign key_original[5274] = key_shuffle[4255];
    assign key_original[5273] = key_shuffle[5572];
    assign key_original[5272] = key_shuffle[5213];
    assign key_original[5271] = key_shuffle[4341];
    assign key_original[5270] = key_shuffle[5000];
    assign key_original[5269] = key_shuffle[4585];
    assign key_original[5268] = key_shuffle[5055];
    assign key_original[5267] = key_shuffle[3775];
    assign key_original[5266] = key_shuffle[6477];
    assign key_original[5265] = key_shuffle[4462];
    assign key_original[5264] = key_shuffle[975];
    assign key_original[5263] = key_shuffle[1712];
    assign key_original[5262] = key_shuffle[7032];
    assign key_original[5261] = key_shuffle[3577];
    assign key_original[5260] = key_shuffle[3984];
    assign key_original[5259] = key_shuffle[3911];
    assign key_original[5258] = key_shuffle[511];
    assign key_original[5257] = key_shuffle[3425];
    assign key_original[5256] = key_shuffle[5338];
    assign key_original[5255] = key_shuffle[5437];
    assign key_original[5254] = key_shuffle[7245];
    assign key_original[5253] = key_shuffle[2594];
    assign key_original[5252] = key_shuffle[2106];
    assign key_original[5251] = key_shuffle[7065];
    assign key_original[5250] = key_shuffle[1686];
    assign key_original[5249] = key_shuffle[668];
    assign key_original[5248] = key_shuffle[932];
    assign key_original[5247] = key_shuffle[613];
    assign key_original[5246] = key_shuffle[4179];
    assign key_original[5245] = key_shuffle[6777];
    assign key_original[5244] = key_shuffle[4634];
    assign key_original[5243] = key_shuffle[4596];
    assign key_original[5242] = key_shuffle[4247];
    assign key_original[5241] = key_shuffle[3369];
    assign key_original[5240] = key_shuffle[7447];
    assign key_original[5239] = key_shuffle[1023];
    assign key_original[5238] = key_shuffle[904];
    assign key_original[5237] = key_shuffle[1876];
    assign key_original[5236] = key_shuffle[3479];
    assign key_original[5235] = key_shuffle[1079];
    assign key_original[5234] = key_shuffle[2316];
    assign key_original[5233] = key_shuffle[117];
    assign key_original[5232] = key_shuffle[945];
    assign key_original[5231] = key_shuffle[296];
    assign key_original[5230] = key_shuffle[5098];
    assign key_original[5229] = key_shuffle[2381];
    assign key_original[5228] = key_shuffle[709];
    assign key_original[5227] = key_shuffle[1302];
    assign key_original[5226] = key_shuffle[7586];
    assign key_original[5225] = key_shuffle[1639];
    assign key_original[5224] = key_shuffle[1287];
    assign key_original[5223] = key_shuffle[3186];
    assign key_original[5222] = key_shuffle[2088];
    assign key_original[5221] = key_shuffle[3061];
    assign key_original[5220] = key_shuffle[937];
    assign key_original[5219] = key_shuffle[1032];
    assign key_original[5218] = key_shuffle[4598];
    assign key_original[5217] = key_shuffle[3599];
    assign key_original[5216] = key_shuffle[4655];
    assign key_original[5215] = key_shuffle[206];
    assign key_original[5214] = key_shuffle[3628];
    assign key_original[5213] = key_shuffle[8069];
    assign key_original[5212] = key_shuffle[7377];
    assign key_original[5211] = key_shuffle[8035];
    assign key_original[5210] = key_shuffle[1471];
    assign key_original[5209] = key_shuffle[6652];
    assign key_original[5208] = key_shuffle[3253];
    assign key_original[5207] = key_shuffle[4727];
    assign key_original[5206] = key_shuffle[1169];
    assign key_original[5205] = key_shuffle[4741];
    assign key_original[5204] = key_shuffle[3653];
    assign key_original[5203] = key_shuffle[6136];
    assign key_original[5202] = key_shuffle[7942];
    assign key_original[5201] = key_shuffle[3810];
    assign key_original[5200] = key_shuffle[1918];
    assign key_original[5199] = key_shuffle[5506];
    assign key_original[5198] = key_shuffle[3231];
    assign key_original[5197] = key_shuffle[4456];
    assign key_original[5196] = key_shuffle[1037];
    assign key_original[5195] = key_shuffle[4821];
    assign key_original[5194] = key_shuffle[2255];
    assign key_original[5193] = key_shuffle[5013];
    assign key_original[5192] = key_shuffle[7530];
    assign key_original[5191] = key_shuffle[6084];
    assign key_original[5190] = key_shuffle[4777];
    assign key_original[5189] = key_shuffle[1518];
    assign key_original[5188] = key_shuffle[4729];
    assign key_original[5187] = key_shuffle[230];
    assign key_original[5186] = key_shuffle[3327];
    assign key_original[5185] = key_shuffle[2590];
    assign key_original[5184] = key_shuffle[5543];
    assign key_original[5183] = key_shuffle[5500];
    assign key_original[5182] = key_shuffle[7008];
    assign key_original[5181] = key_shuffle[983];
    assign key_original[5180] = key_shuffle[3418];
    assign key_original[5179] = key_shuffle[3004];
    assign key_original[5178] = key_shuffle[6014];
    assign key_original[5177] = key_shuffle[3794];
    assign key_original[5176] = key_shuffle[1433];
    assign key_original[5175] = key_shuffle[2017];
    assign key_original[5174] = key_shuffle[6922];
    assign key_original[5173] = key_shuffle[4282];
    assign key_original[5172] = key_shuffle[7497];
    assign key_original[5171] = key_shuffle[7928];
    assign key_original[5170] = key_shuffle[6246];
    assign key_original[5169] = key_shuffle[7316];
    assign key_original[5168] = key_shuffle[5526];
    assign key_original[5167] = key_shuffle[4626];
    assign key_original[5166] = key_shuffle[4416];
    assign key_original[5165] = key_shuffle[2894];
    assign key_original[5164] = key_shuffle[6288];
    assign key_original[5163] = key_shuffle[3134];
    assign key_original[5162] = key_shuffle[5340];
    assign key_original[5161] = key_shuffle[3933];
    assign key_original[5160] = key_shuffle[1087];
    assign key_original[5159] = key_shuffle[3388];
    assign key_original[5158] = key_shuffle[6516];
    assign key_original[5157] = key_shuffle[3089];
    assign key_original[5156] = key_shuffle[2109];
    assign key_original[5155] = key_shuffle[4133];
    assign key_original[5154] = key_shuffle[2642];
    assign key_original[5153] = key_shuffle[6565];
    assign key_original[5152] = key_shuffle[4611];
    assign key_original[5151] = key_shuffle[2156];
    assign key_original[5150] = key_shuffle[1268];
    assign key_original[5149] = key_shuffle[3630];
    assign key_original[5148] = key_shuffle[2482];
    assign key_original[5147] = key_shuffle[6676];
    assign key_original[5146] = key_shuffle[2569];
    assign key_original[5145] = key_shuffle[5870];
    assign key_original[5144] = key_shuffle[4804];
    assign key_original[5143] = key_shuffle[7039];
    assign key_original[5142] = key_shuffle[334];
    assign key_original[5141] = key_shuffle[1059];
    assign key_original[5140] = key_shuffle[4427];
    assign key_original[5139] = key_shuffle[6468];
    assign key_original[5138] = key_shuffle[2401];
    assign key_original[5137] = key_shuffle[2965];
    assign key_original[5136] = key_shuffle[4935];
    assign key_original[5135] = key_shuffle[214];
    assign key_original[5134] = key_shuffle[3276];
    assign key_original[5133] = key_shuffle[4285];
    assign key_original[5132] = key_shuffle[4372];
    assign key_original[5131] = key_shuffle[3021];
    assign key_original[5130] = key_shuffle[3865];
    assign key_original[5129] = key_shuffle[3398];
    assign key_original[5128] = key_shuffle[5419];
    assign key_original[5127] = key_shuffle[6397];
    assign key_original[5126] = key_shuffle[1303];
    assign key_original[5125] = key_shuffle[6843];
    assign key_original[5124] = key_shuffle[228];
    assign key_original[5123] = key_shuffle[2391];
    assign key_original[5122] = key_shuffle[6649];
    assign key_original[5121] = key_shuffle[2787];
    assign key_original[5120] = key_shuffle[4033];
    assign key_original[5119] = key_shuffle[4248];
    assign key_original[5118] = key_shuffle[4815];
    assign key_original[5117] = key_shuffle[7663];
    assign key_original[5116] = key_shuffle[4328];
    assign key_original[5115] = key_shuffle[6248];
    assign key_original[5114] = key_shuffle[2030];
    assign key_original[5113] = key_shuffle[4195];
    assign key_original[5112] = key_shuffle[833];
    assign key_original[5111] = key_shuffle[1540];
    assign key_original[5110] = key_shuffle[1728];
    assign key_original[5109] = key_shuffle[6364];
    assign key_original[5108] = key_shuffle[2034];
    assign key_original[5107] = key_shuffle[3447];
    assign key_original[5106] = key_shuffle[3528];
    assign key_original[5105] = key_shuffle[1726];
    assign key_original[5104] = key_shuffle[2818];
    assign key_original[5103] = key_shuffle[7861];
    assign key_original[5102] = key_shuffle[3050];
    assign key_original[5101] = key_shuffle[7617];
    assign key_original[5100] = key_shuffle[743];
    assign key_original[5099] = key_shuffle[2954];
    assign key_original[5098] = key_shuffle[3386];
    assign key_original[5097] = key_shuffle[7212];
    assign key_original[5096] = key_shuffle[2842];
    assign key_original[5095] = key_shuffle[5619];
    assign key_original[5094] = key_shuffle[964];
    assign key_original[5093] = key_shuffle[1470];
    assign key_original[5092] = key_shuffle[788];
    assign key_original[5091] = key_shuffle[1602];
    assign key_original[5090] = key_shuffle[3318];
    assign key_original[5089] = key_shuffle[5481];
    assign key_original[5088] = key_shuffle[1236];
    assign key_original[5087] = key_shuffle[3961];
    assign key_original[5086] = key_shuffle[7100];
    assign key_original[5085] = key_shuffle[6205];
    assign key_original[5084] = key_shuffle[2596];
    assign key_original[5083] = key_shuffle[635];
    assign key_original[5082] = key_shuffle[6219];
    assign key_original[5081] = key_shuffle[2179];
    assign key_original[5080] = key_shuffle[5347];
    assign key_original[5079] = key_shuffle[796];
    assign key_original[5078] = key_shuffle[7895];
    assign key_original[5077] = key_shuffle[7287];
    assign key_original[5076] = key_shuffle[7544];
    assign key_original[5075] = key_shuffle[5420];
    assign key_original[5074] = key_shuffle[4464];
    assign key_original[5073] = key_shuffle[4007];
    assign key_original[5072] = key_shuffle[5431];
    assign key_original[5071] = key_shuffle[6194];
    assign key_original[5070] = key_shuffle[5175];
    assign key_original[5069] = key_shuffle[5067];
    assign key_original[5068] = key_shuffle[2575];
    assign key_original[5067] = key_shuffle[2365];
    assign key_original[5066] = key_shuffle[175];
    assign key_original[5065] = key_shuffle[6532];
    assign key_original[5064] = key_shuffle[380];
    assign key_original[5063] = key_shuffle[5111];
    assign key_original[5062] = key_shuffle[8096];
    assign key_original[5061] = key_shuffle[6590];
    assign key_original[5060] = key_shuffle[3091];
    assign key_original[5059] = key_shuffle[3953];
    assign key_original[5058] = key_shuffle[5843];
    assign key_original[5057] = key_shuffle[7290];
    assign key_original[5056] = key_shuffle[3185];
    assign key_original[5055] = key_shuffle[7609];
    assign key_original[5054] = key_shuffle[2501];
    assign key_original[5053] = key_shuffle[3483];
    assign key_original[5052] = key_shuffle[1968];
    assign key_original[5051] = key_shuffle[8113];
    assign key_original[5050] = key_shuffle[7956];
    assign key_original[5049] = key_shuffle[3103];
    assign key_original[5048] = key_shuffle[7997];
    assign key_original[5047] = key_shuffle[3951];
    assign key_original[5046] = key_shuffle[577];
    assign key_original[5045] = key_shuffle[6631];
    assign key_original[5044] = key_shuffle[4619];
    assign key_original[5043] = key_shuffle[4948];
    assign key_original[5042] = key_shuffle[1981];
    assign key_original[5041] = key_shuffle[5007];
    assign key_original[5040] = key_shuffle[5835];
    assign key_original[5039] = key_shuffle[2717];
    assign key_original[5038] = key_shuffle[1758];
    assign key_original[5037] = key_shuffle[4449];
    assign key_original[5036] = key_shuffle[959];
    assign key_original[5035] = key_shuffle[5010];
    assign key_original[5034] = key_shuffle[2007];
    assign key_original[5033] = key_shuffle[6471];
    assign key_original[5032] = key_shuffle[1811];
    assign key_original[5031] = key_shuffle[4024];
    assign key_original[5030] = key_shuffle[4601];
    assign key_original[5029] = key_shuffle[4569];
    assign key_original[5028] = key_shuffle[2437];
    assign key_original[5027] = key_shuffle[5287];
    assign key_original[5026] = key_shuffle[6332];
    assign key_original[5025] = key_shuffle[7994];
    assign key_original[5024] = key_shuffle[6604];
    assign key_original[5023] = key_shuffle[3412];
    assign key_original[5022] = key_shuffle[7794];
    assign key_original[5021] = key_shuffle[2653];
    assign key_original[5020] = key_shuffle[5259];
    assign key_original[5019] = key_shuffle[7342];
    assign key_original[5018] = key_shuffle[6946];
    assign key_original[5017] = key_shuffle[2303];
    assign key_original[5016] = key_shuffle[6166];
    assign key_original[5015] = key_shuffle[4771];
    assign key_original[5014] = key_shuffle[1907];
    assign key_original[5013] = key_shuffle[4961];
    assign key_original[5012] = key_shuffle[3331];
    assign key_original[5011] = key_shuffle[4223];
    assign key_original[5010] = key_shuffle[3079];
    assign key_original[5009] = key_shuffle[398];
    assign key_original[5008] = key_shuffle[5573];
    assign key_original[5007] = key_shuffle[6690];
    assign key_original[5006] = key_shuffle[3219];
    assign key_original[5005] = key_shuffle[1036];
    assign key_original[5004] = key_shuffle[4938];
    assign key_original[5003] = key_shuffle[1006];
    assign key_original[5002] = key_shuffle[6759];
    assign key_original[5001] = key_shuffle[761];
    assign key_original[5000] = key_shuffle[378];
    assign key_original[4999] = key_shuffle[7321];
    assign key_original[4998] = key_shuffle[129];
    assign key_original[4997] = key_shuffle[4076];
    assign key_original[4996] = key_shuffle[1056];
    assign key_original[4995] = key_shuffle[1209];
    assign key_original[4994] = key_shuffle[7587];
    assign key_original[4993] = key_shuffle[2172];
    assign key_original[4992] = key_shuffle[6167];
    assign key_original[4991] = key_shuffle[490];
    assign key_original[4990] = key_shuffle[974];
    assign key_original[4989] = key_shuffle[4051];
    assign key_original[4988] = key_shuffle[3169];
    assign key_original[4987] = key_shuffle[2705];
    assign key_original[4986] = key_shuffle[6000];
    assign key_original[4985] = key_shuffle[3645];
    assign key_original[4984] = key_shuffle[5295];
    assign key_original[4983] = key_shuffle[4453];
    assign key_original[4982] = key_shuffle[7387];
    assign key_original[4981] = key_shuffle[3178];
    assign key_original[4980] = key_shuffle[1045];
    assign key_original[4979] = key_shuffle[3756];
    assign key_original[4978] = key_shuffle[4990];
    assign key_original[4977] = key_shuffle[1485];
    assign key_original[4976] = key_shuffle[4316];
    assign key_original[4975] = key_shuffle[6199];
    assign key_original[4974] = key_shuffle[8124];
    assign key_original[4973] = key_shuffle[1458];
    assign key_original[4972] = key_shuffle[1722];
    assign key_original[4971] = key_shuffle[8055];
    assign key_original[4970] = key_shuffle[7104];
    assign key_original[4969] = key_shuffle[4923];
    assign key_original[4968] = key_shuffle[6176];
    assign key_original[4967] = key_shuffle[6818];
    assign key_original[4966] = key_shuffle[1685];
    assign key_original[4965] = key_shuffle[2755];
    assign key_original[4964] = key_shuffle[159];
    assign key_original[4963] = key_shuffle[3815];
    assign key_original[4962] = key_shuffle[7723];
    assign key_original[4961] = key_shuffle[5048];
    assign key_original[4960] = key_shuffle[5240];
    assign key_original[4959] = key_shuffle[1389];
    assign key_original[4958] = key_shuffle[3419];
    assign key_original[4957] = key_shuffle[6842];
    assign key_original[4956] = key_shuffle[6131];
    assign key_original[4955] = key_shuffle[3633];
    assign key_original[4954] = key_shuffle[5265];
    assign key_original[4953] = key_shuffle[2229];
    assign key_original[4952] = key_shuffle[644];
    assign key_original[4951] = key_shuffle[1380];
    assign key_original[4950] = key_shuffle[8016];
    assign key_original[4949] = key_shuffle[2282];
    assign key_original[4948] = key_shuffle[3861];
    assign key_original[4947] = key_shuffle[5170];
    assign key_original[4946] = key_shuffle[5525];
    assign key_original[4945] = key_shuffle[4883];
    assign key_original[4944] = key_shuffle[8176];
    assign key_original[4943] = key_shuffle[4376];
    assign key_original[4942] = key_shuffle[39];
    assign key_original[4941] = key_shuffle[4260];
    assign key_original[4940] = key_shuffle[7882];
    assign key_original[4939] = key_shuffle[6201];
    assign key_original[4938] = key_shuffle[472];
    assign key_original[4937] = key_shuffle[3921];
    assign key_original[4936] = key_shuffle[3151];
    assign key_original[4935] = key_shuffle[8057];
    assign key_original[4934] = key_shuffle[809];
    assign key_original[4933] = key_shuffle[1359];
    assign key_original[4932] = key_shuffle[1710];
    assign key_original[4931] = key_shuffle[5196];
    assign key_original[4930] = key_shuffle[2587];
    assign key_original[4929] = key_shuffle[5827];
    assign key_original[4928] = key_shuffle[2238];
    assign key_original[4927] = key_shuffle[1891];
    assign key_original[4926] = key_shuffle[2966];
    assign key_original[4925] = key_shuffle[6855];
    assign key_original[4924] = key_shuffle[4653];
    assign key_original[4923] = key_shuffle[4040];
    assign key_original[4922] = key_shuffle[6299];
    assign key_original[4921] = key_shuffle[5885];
    assign key_original[4920] = key_shuffle[7759];
    assign key_original[4919] = key_shuffle[1729];
    assign key_original[4918] = key_shuffle[5529];
    assign key_original[4917] = key_shuffle[7003];
    assign key_original[4916] = key_shuffle[1893];
    assign key_original[4915] = key_shuffle[4230];
    assign key_original[4914] = key_shuffle[7533];
    assign key_original[4913] = key_shuffle[7439];
    assign key_original[4912] = key_shuffle[3855];
    assign key_original[4911] = key_shuffle[6748];
    assign key_original[4910] = key_shuffle[1829];
    assign key_original[4909] = key_shuffle[6203];
    assign key_original[4908] = key_shuffle[2173];
    assign key_original[4907] = key_shuffle[7705];
    assign key_original[4906] = key_shuffle[3022];
    assign key_original[4905] = key_shuffle[2470];
    assign key_original[4904] = key_shuffle[6605];
    assign key_original[4903] = key_shuffle[6300];
    assign key_original[4902] = key_shuffle[7970];
    assign key_original[4901] = key_shuffle[7186];
    assign key_original[4900] = key_shuffle[1506];
    assign key_original[4899] = key_shuffle[5975];
    assign key_original[4898] = key_shuffle[250];
    assign key_original[4897] = key_shuffle[7315];
    assign key_original[4896] = key_shuffle[6802];
    assign key_original[4895] = key_shuffle[3862];
    assign key_original[4894] = key_shuffle[6452];
    assign key_original[4893] = key_shuffle[6766];
    assign key_original[4892] = key_shuffle[721];
    assign key_original[4891] = key_shuffle[7128];
    assign key_original[4890] = key_shuffle[1814];
    assign key_original[4889] = key_shuffle[7616];
    assign key_original[4888] = key_shuffle[144];
    assign key_original[4887] = key_shuffle[1128];
    assign key_original[4886] = key_shuffle[6382];
    assign key_original[4885] = key_shuffle[4043];
    assign key_original[4884] = key_shuffle[1158];
    assign key_original[4883] = key_shuffle[6261];
    assign key_original[4882] = key_shuffle[279];
    assign key_original[4881] = key_shuffle[7519];
    assign key_original[4880] = key_shuffle[238];
    assign key_original[4879] = key_shuffle[7108];
    assign key_original[4878] = key_shuffle[5315];
    assign key_original[4877] = key_shuffle[3391];
    assign key_original[4876] = key_shuffle[7449];
    assign key_original[4875] = key_shuffle[2163];
    assign key_original[4874] = key_shuffle[4915];
    assign key_original[4873] = key_shuffle[7792];
    assign key_original[4872] = key_shuffle[7789];
    assign key_original[4871] = key_shuffle[2861];
    assign key_original[4870] = key_shuffle[1711];
    assign key_original[4869] = key_shuffle[2148];
    assign key_original[4868] = key_shuffle[5880];
    assign key_original[4867] = key_shuffle[4369];
    assign key_original[4866] = key_shuffle[2836];
    assign key_original[4865] = key_shuffle[1886];
    assign key_original[4864] = key_shuffle[2519];
    assign key_original[4863] = key_shuffle[164];
    assign key_original[4862] = key_shuffle[3787];
    assign key_original[4861] = key_shuffle[1837];
    assign key_original[4860] = key_shuffle[370];
    assign key_original[4859] = key_shuffle[6755];
    assign key_original[4858] = key_shuffle[741];
    assign key_original[4857] = key_shuffle[5412];
    assign key_original[4856] = key_shuffle[1642];
    assign key_original[4855] = key_shuffle[4045];
    assign key_original[4854] = key_shuffle[5220];
    assign key_original[4853] = key_shuffle[7219];
    assign key_original[4852] = key_shuffle[26];
    assign key_original[4851] = key_shuffle[512];
    assign key_original[4850] = key_shuffle[2064];
    assign key_original[4849] = key_shuffle[5736];
    assign key_original[4848] = key_shuffle[2908];
    assign key_original[4847] = key_shuffle[3902];
    assign key_original[4846] = key_shuffle[5074];
    assign key_original[4845] = key_shuffle[1664];
    assign key_original[4844] = key_shuffle[6744];
    assign key_original[4843] = key_shuffle[5509];
    assign key_original[4842] = key_shuffle[3212];
    assign key_original[4841] = key_shuffle[358];
    assign key_original[4840] = key_shuffle[6075];
    assign key_original[4839] = key_shuffle[2855];
    assign key_original[4838] = key_shuffle[1203];
    assign key_original[4837] = key_shuffle[4252];
    assign key_original[4836] = key_shuffle[4739];
    assign key_original[4835] = key_shuffle[7930];
    assign key_original[4834] = key_shuffle[2976];
    assign key_original[4833] = key_shuffle[1670];
    assign key_original[4832] = key_shuffle[6753];
    assign key_original[4831] = key_shuffle[5779];
    assign key_original[4830] = key_shuffle[7107];
    assign key_original[4829] = key_shuffle[2253];
    assign key_original[4828] = key_shuffle[6756];
    assign key_original[4827] = key_shuffle[2631];
    assign key_original[4826] = key_shuffle[2359];
    assign key_original[4825] = key_shuffle[141];
    assign key_original[4824] = key_shuffle[1553];
    assign key_original[4823] = key_shuffle[2374];
    assign key_original[4822] = key_shuffle[5254];
    assign key_original[4821] = key_shuffle[553];
    assign key_original[4820] = key_shuffle[6407];
    assign key_original[4819] = key_shuffle[7624];
    assign key_original[4818] = key_shuffle[4295];
    assign key_original[4817] = key_shuffle[877];
    assign key_original[4816] = key_shuffle[4269];
    assign key_original[4815] = key_shuffle[4074];
    assign key_original[4814] = key_shuffle[3395];
    assign key_original[4813] = key_shuffle[7976];
    assign key_original[4812] = key_shuffle[1716];
    assign key_original[4811] = key_shuffle[655];
    assign key_original[4810] = key_shuffle[353];
    assign key_original[4809] = key_shuffle[7579];
    assign key_original[4808] = key_shuffle[1815];
    assign key_original[4807] = key_shuffle[1142];
    assign key_original[4806] = key_shuffle[3394];
    assign key_original[4805] = key_shuffle[4870];
    assign key_original[4804] = key_shuffle[1597];
    assign key_original[4803] = key_shuffle[2700];
    assign key_original[4802] = key_shuffle[17];
    assign key_original[4801] = key_shuffle[715];
    assign key_original[4800] = key_shuffle[5981];
    assign key_original[4799] = key_shuffle[3148];
    assign key_original[4798] = key_shuffle[3590];
    assign key_original[4797] = key_shuffle[5681];
    assign key_original[4796] = key_shuffle[3161];
    assign key_original[4795] = key_shuffle[6331];
    assign key_original[4794] = key_shuffle[7751];
    assign key_original[4793] = key_shuffle[1509];
    assign key_original[4792] = key_shuffle[3644];
    assign key_original[4791] = key_shuffle[6037];
    assign key_original[4790] = key_shuffle[4406];
    assign key_original[4789] = key_shuffle[6513];
    assign key_original[4788] = key_shuffle[1966];
    assign key_original[4787] = key_shuffle[4681];
    assign key_original[4786] = key_shuffle[7729];
    assign key_original[4785] = key_shuffle[426];
    assign key_original[4784] = key_shuffle[4884];
    assign key_original[4783] = key_shuffle[3462];
    assign key_original[4782] = key_shuffle[6677];
    assign key_original[4781] = key_shuffle[2986];
    assign key_original[4780] = key_shuffle[2318];
    assign key_original[4779] = key_shuffle[7721];
    assign key_original[4778] = key_shuffle[915];
    assign key_original[4777] = key_shuffle[1035];
    assign key_original[4776] = key_shuffle[1365];
    assign key_original[4775] = key_shuffle[768];
    assign key_original[4774] = key_shuffle[6209];
    assign key_original[4773] = key_shuffle[5855];
    assign key_original[4772] = key_shuffle[2290];
    assign key_original[4771] = key_shuffle[1192];
    assign key_original[4770] = key_shuffle[7283];
    assign key_original[4769] = key_shuffle[7604];
    assign key_original[4768] = key_shuffle[6783];
    assign key_original[4767] = key_shuffle[375];
    assign key_original[4766] = key_shuffle[2310];
    assign key_original[4765] = key_shuffle[6616];
    assign key_original[4764] = key_shuffle[6294];
    assign key_original[4763] = key_shuffle[2781];
    assign key_original[4762] = key_shuffle[5618];
    assign key_original[4761] = key_shuffle[5657];
    assign key_original[4760] = key_shuffle[1333];
    assign key_original[4759] = key_shuffle[3635];
    assign key_original[4758] = key_shuffle[7554];
    assign key_original[4757] = key_shuffle[327];
    assign key_original[4756] = key_shuffle[820];
    assign key_original[4755] = key_shuffle[5992];
    assign key_original[4754] = key_shuffle[6048];
    assign key_original[4753] = key_shuffle[2424];
    assign key_original[4752] = key_shuffle[3832];
    assign key_original[4751] = key_shuffle[1388];
    assign key_original[4750] = key_shuffle[5560];
    assign key_original[4749] = key_shuffle[2458];
    assign key_original[4748] = key_shuffle[5330];
    assign key_original[4747] = key_shuffle[4861];
    assign key_original[4746] = key_shuffle[2048];
    assign key_original[4745] = key_shuffle[7815];
    assign key_original[4744] = key_shuffle[5408];
    assign key_original[4743] = key_shuffle[2296];
    assign key_original[4742] = key_shuffle[6850];
    assign key_original[4741] = key_shuffle[7299];
    assign key_original[4740] = key_shuffle[1223];
    assign key_original[4739] = key_shuffle[229];
    assign key_original[4738] = key_shuffle[3602];
    assign key_original[4737] = key_shuffle[5263];
    assign key_original[4736] = key_shuffle[6025];
    assign key_original[4735] = key_shuffle[5632];
    assign key_original[4734] = key_shuffle[6600];
    assign key_original[4733] = key_shuffle[1961];
    assign key_original[4732] = key_shuffle[4776];
    assign key_original[4731] = key_shuffle[783];
    assign key_original[4730] = key_shuffle[4366];
    assign key_original[4729] = key_shuffle[2579];
    assign key_original[4728] = key_shuffle[2160];
    assign key_original[4727] = key_shuffle[657];
    assign key_original[4726] = key_shuffle[520];
    assign key_original[4725] = key_shuffle[4335];
    assign key_original[4724] = key_shuffle[6546];
    assign key_original[4723] = key_shuffle[4420];
    assign key_original[4722] = key_shuffle[6465];
    assign key_original[4721] = key_shuffle[6933];
    assign key_original[4720] = key_shuffle[3739];
    assign key_original[4719] = key_shuffle[7084];
    assign key_original[4718] = key_shuffle[1420];
    assign key_original[4717] = key_shuffle[4885];
    assign key_original[4716] = key_shuffle[1304];
    assign key_original[4715] = key_shuffle[962];
    assign key_original[4714] = key_shuffle[722];
    assign key_original[4713] = key_shuffle[2323];
    assign key_original[4712] = key_shuffle[8157];
    assign key_original[4711] = key_shuffle[5866];
    assign key_original[4710] = key_shuffle[163];
    assign key_original[4709] = key_shuffle[2820];
    assign key_original[4708] = key_shuffle[6702];
    assign key_original[4707] = key_shuffle[8008];
    assign key_original[4706] = key_shuffle[6071];
    assign key_original[4705] = key_shuffle[4807];
    assign key_original[4704] = key_shuffle[1884];
    assign key_original[4703] = key_shuffle[797];
    assign key_original[4702] = key_shuffle[7382];
    assign key_original[4701] = key_shuffle[4281];
    assign key_original[4700] = key_shuffle[3107];
    assign key_original[4699] = key_shuffle[112];
    assign key_original[4698] = key_shuffle[271];
    assign key_original[4697] = key_shuffle[106];
    assign key_original[4696] = key_shuffle[1439];
    assign key_original[4695] = key_shuffle[1915];
    assign key_original[4694] = key_shuffle[2526];
    assign key_original[4693] = key_shuffle[4906];
    assign key_original[4692] = key_shuffle[3655];
    assign key_original[4691] = key_shuffle[1355];
    assign key_original[4690] = key_shuffle[6271];
    assign key_original[4689] = key_shuffle[1840];
    assign key_original[4688] = key_shuffle[5757];
    assign key_original[4687] = key_shuffle[2989];
    assign key_original[4686] = key_shuffle[7370];
    assign key_original[4685] = key_shuffle[8009];
    assign key_original[4684] = key_shuffle[6872];
    assign key_original[4683] = key_shuffle[3081];
    assign key_original[4682] = key_shuffle[1587];
    assign key_original[4681] = key_shuffle[4610];
    assign key_original[4680] = key_shuffle[6390];
    assign key_original[4679] = key_shuffle[5394];
    assign key_original[4678] = key_shuffle[4428];
    assign key_original[4677] = key_shuffle[5941];
    assign key_original[4676] = key_shuffle[3244];
    assign key_original[4675] = key_shuffle[270];
    assign key_original[4674] = key_shuffle[5277];
    assign key_original[4673] = key_shuffle[1769];
    assign key_original[4672] = key_shuffle[7465];
    assign key_original[4671] = key_shuffle[7501];
    assign key_original[4670] = key_shuffle[7206];
    assign key_original[4669] = key_shuffle[4351];
    assign key_original[4668] = key_shuffle[2979];
    assign key_original[4667] = key_shuffle[6366];
    assign key_original[4666] = key_shuffle[2293];
    assign key_original[4665] = key_shuffle[7295];
    assign key_original[4664] = key_shuffle[3401];
    assign key_original[4663] = key_shuffle[1663];
    assign key_original[4662] = key_shuffle[1031];
    assign key_original[4661] = key_shuffle[5792];
    assign key_original[4660] = key_shuffle[689];
    assign key_original[4659] = key_shuffle[1372];
    assign key_original[4658] = key_shuffle[1946];
    assign key_original[4657] = key_shuffle[2039];
    assign key_original[4656] = key_shuffle[7653];
    assign key_original[4655] = key_shuffle[6019];
    assign key_original[4654] = key_shuffle[6126];
    assign key_original[4653] = key_shuffle[7004];
    assign key_original[4652] = key_shuffle[4146];
    assign key_original[4651] = key_shuffle[3410];
    assign key_original[4650] = key_shuffle[3748];
    assign key_original[4649] = key_shuffle[5327];
    assign key_original[4648] = key_shuffle[4307];
    assign key_original[4647] = key_shuffle[5291];
    assign key_original[4646] = key_shuffle[794];
    assign key_original[4645] = key_shuffle[3137];
    assign key_original[4644] = key_shuffle[5939];
    assign key_original[4643] = key_shuffle[7854];
    assign key_original[4642] = key_shuffle[6046];
    assign key_original[4641] = key_shuffle[1057];
    assign key_original[4640] = key_shuffle[1395];
    assign key_original[4639] = key_shuffle[4997];
    assign key_original[4638] = key_shuffle[2612];
    assign key_original[4637] = key_shuffle[2184];
    assign key_original[4636] = key_shuffle[5640];
    assign key_original[4635] = key_shuffle[8159];
    assign key_original[4634] = key_shuffle[59];
    assign key_original[4633] = key_shuffle[7062];
    assign key_original[4632] = key_shuffle[3016];
    assign key_original[4631] = key_shuffle[3452];
    assign key_original[4630] = key_shuffle[5977];
    assign key_original[4629] = key_shuffle[3976];
    assign key_original[4628] = key_shuffle[2548];
    assign key_original[4627] = key_shuffle[1900];
    assign key_original[4626] = key_shuffle[7906];
    assign key_original[4625] = key_shuffle[4786];
    assign key_original[4624] = key_shuffle[2123];
    assign key_original[4623] = key_shuffle[2828];
    assign key_original[4622] = key_shuffle[1730];
    assign key_original[4621] = key_shuffle[7612];
    assign key_original[4620] = key_shuffle[3046];
    assign key_original[4619] = key_shuffle[2623];
    assign key_original[4618] = key_shuffle[1522];
    assign key_original[4617] = key_shuffle[2927];
    assign key_original[4616] = key_shuffle[4434];
    assign key_original[4615] = key_shuffle[5432];
    assign key_original[4614] = key_shuffle[342];
    assign key_original[4613] = key_shuffle[1611];
    assign key_original[4612] = key_shuffle[7293];
    assign key_original[4611] = key_shuffle[6247];
    assign key_original[4610] = key_shuffle[2739];
    assign key_original[4609] = key_shuffle[4149];
    assign key_original[4608] = key_shuffle[2295];
    assign key_original[4607] = key_shuffle[7784];
    assign key_original[4606] = key_shuffle[587];
    assign key_original[4605] = key_shuffle[776];
    assign key_original[4604] = key_shuffle[3626];
    assign key_original[4603] = key_shuffle[1654];
    assign key_original[4602] = key_shuffle[5378];
    assign key_original[4601] = key_shuffle[5630];
    assign key_original[4600] = key_shuffle[3508];
    assign key_original[4599] = key_shuffle[4280];
    assign key_original[4598] = key_shuffle[1460];
    assign key_original[4597] = key_shuffle[4738];
    assign key_original[4596] = key_shuffle[468];
    assign key_original[4595] = key_shuffle[7915];
    assign key_original[4594] = key_shuffle[3157];
    assign key_original[4593] = key_shuffle[7095];
    assign key_original[4592] = key_shuffle[3007];
    assign key_original[4591] = key_shuffle[6442];
    assign key_original[4590] = key_shuffle[3190];
    assign key_original[4589] = key_shuffle[6960];
    assign key_original[4588] = key_shuffle[5717];
    assign key_original[4587] = key_shuffle[1277];
    assign key_original[4586] = key_shuffle[3380];
    assign key_original[4585] = key_shuffle[7049];
    assign key_original[4584] = key_shuffle[6899];
    assign key_original[4583] = key_shuffle[884];
    assign key_original[4582] = key_shuffle[5728];
    assign key_original[4581] = key_shuffle[2399];
    assign key_original[4580] = key_shuffle[1610];
    assign key_original[4579] = key_shuffle[6385];
    assign key_original[4578] = key_shuffle[38];
    assign key_original[4577] = key_shuffle[515];
    assign key_original[4576] = key_shuffle[6374];
    assign key_original[4575] = key_shuffle[1619];
    assign key_original[4574] = key_shuffle[2841];
    assign key_original[4573] = key_shuffle[5721];
    assign key_original[4572] = key_shuffle[7774];
    assign key_original[4571] = key_shuffle[389];
    assign key_original[4570] = key_shuffle[2628];
    assign key_original[4569] = key_shuffle[2009];
    assign key_original[4568] = key_shuffle[5893];
    assign key_original[4567] = key_shuffle[4993];
    assign key_original[4566] = key_shuffle[4828];
    assign key_original[4565] = key_shuffle[1296];
    assign key_original[4564] = key_shuffle[3272];
    assign key_original[4563] = key_shuffle[3135];
    assign key_original[4562] = key_shuffle[4436];
    assign key_original[4561] = key_shuffle[1472];
    assign key_original[4560] = key_shuffle[5363];
    assign key_original[4559] = key_shuffle[1860];
    assign key_original[4558] = key_shuffle[602];
    assign key_original[4557] = key_shuffle[2085];
    assign key_original[4556] = key_shuffle[984];
    assign key_original[4555] = key_shuffle[170];
    assign key_original[4554] = key_shuffle[3947];
    assign key_original[4553] = key_shuffle[6651];
    assign key_original[4552] = key_shuffle[6425];
    assign key_original[4551] = key_shuffle[967];
    assign key_original[4550] = key_shuffle[7199];
    assign key_original[4549] = key_shuffle[1909];
    assign key_original[4548] = key_shuffle[1844];
    assign key_original[4547] = key_shuffle[1958];
    assign key_original[4546] = key_shuffle[6123];
    assign key_original[4545] = key_shuffle[1384];
    assign key_original[4544] = key_shuffle[3588];
    assign key_original[4543] = key_shuffle[4017];
    assign key_original[4542] = key_shuffle[4812];
    assign key_original[4541] = key_shuffle[3225];
    assign key_original[4540] = key_shuffle[4233];
    assign key_original[4539] = key_shuffle[1094];
    assign key_original[4538] = key_shuffle[4896];
    assign key_original[4537] = key_shuffle[7075];
    assign key_original[4536] = key_shuffle[7090];
    assign key_original[4535] = key_shuffle[2161];
    assign key_original[4534] = key_shuffle[3220];
    assign key_original[4533] = key_shuffle[7374];
    assign key_original[4532] = key_shuffle[7088];
    assign key_original[4531] = key_shuffle[2093];
    assign key_original[4530] = key_shuffle[1974];
    assign key_original[4529] = key_shuffle[2649];
    assign key_original[4528] = key_shuffle[3048];
    assign key_original[4527] = key_shuffle[2199];
    assign key_original[4526] = key_shuffle[2393];
    assign key_original[4525] = key_shuffle[2538];
    assign key_original[4524] = key_shuffle[7052];
    assign key_original[4523] = key_shuffle[760];
    assign key_original[4522] = key_shuffle[2663];
    assign key_original[4521] = key_shuffle[1740];
    assign key_original[4520] = key_shuffle[532];
    assign key_original[4519] = key_shuffle[7829];
    assign key_original[4518] = key_shuffle[1456];
    assign key_original[4517] = key_shuffle[7570];
    assign key_original[4516] = key_shuffle[5921];
    assign key_original[4515] = key_shuffle[2912];
    assign key_original[4514] = key_shuffle[664];
    assign key_original[4513] = key_shuffle[4740];
    assign key_original[4512] = key_shuffle[138];
    assign key_original[4511] = key_shuffle[7949];
    assign key_original[4510] = key_shuffle[83];
    assign key_original[4509] = key_shuffle[7989];
    assign key_original[4508] = key_shuffle[3040];
    assign key_original[4507] = key_shuffle[6852];
    assign key_original[4506] = key_shuffle[7269];
    assign key_original[4505] = key_shuffle[539];
    assign key_original[4504] = key_shuffle[414];
    assign key_original[4503] = key_shuffle[7426];
    assign key_original[4502] = key_shuffle[3687];
    assign key_original[4501] = key_shuffle[4921];
    assign key_original[4500] = key_shuffle[3130];
    assign key_original[4499] = key_shuffle[6021];
    assign key_original[4498] = key_shuffle[2956];
    assign key_original[4497] = key_shuffle[3703];
    assign key_original[4496] = key_shuffle[2278];
    assign key_original[4495] = key_shuffle[162];
    assign key_original[4494] = key_shuffle[5689];
    assign key_original[4493] = key_shuffle[1749];
    assign key_original[4492] = key_shuffle[6542];
    assign key_original[4491] = key_shuffle[1483];
    assign key_original[4490] = key_shuffle[5650];
    assign key_original[4489] = key_shuffle[2611];
    assign key_original[4488] = key_shuffle[5480];
    assign key_original[4487] = key_shuffle[1077];
    assign key_original[4486] = key_shuffle[1906];
    assign key_original[4485] = key_shuffle[4696];
    assign key_original[4484] = key_shuffle[7712];
    assign key_original[4483] = key_shuffle[6624];
    assign key_original[4482] = key_shuffle[427];
    assign key_original[4481] = key_shuffle[4617];
    assign key_original[4480] = key_shuffle[5056];
    assign key_original[4479] = key_shuffle[3847];
    assign key_original[4478] = key_shuffle[4240];
    assign key_original[4477] = key_shuffle[3586];
    assign key_original[4476] = key_shuffle[7495];
    assign key_original[4475] = key_shuffle[1489];
    assign key_original[4474] = key_shuffle[5211];
    assign key_original[4473] = key_shuffle[943];
    assign key_original[4472] = key_shuffle[1615];
    assign key_original[4471] = key_shuffle[3881];
    assign key_original[4470] = key_shuffle[2536];
    assign key_original[4469] = key_shuffle[4030];
    assign key_original[4468] = key_shuffle[6586];
    assign key_original[4467] = key_shuffle[5963];
    assign key_original[4466] = key_shuffle[6121];
    assign key_original[4465] = key_shuffle[3542];
    assign key_original[4464] = key_shuffle[7818];
    assign key_original[4463] = key_shuffle[5710];
    assign key_original[4462] = key_shuffle[764];
    assign key_original[4461] = key_shuffle[6128];
    assign key_original[4460] = key_shuffle[7129];
    assign key_original[4459] = key_shuffle[4209];
    assign key_original[4458] = key_shuffle[78];
    assign key_original[4457] = key_shuffle[4743];
    assign key_original[4456] = key_shuffle[1865];
    assign key_original[4455] = key_shuffle[503];
    assign key_original[4454] = key_shuffle[3662];
    assign key_original[4453] = key_shuffle[1924];
    assign key_original[4452] = key_shuffle[5197];
    assign key_original[4451] = key_shuffle[2751];
    assign key_original[4450] = key_shuffle[970];
    assign key_original[4449] = key_shuffle[2089];
    assign key_original[4448] = key_shuffle[7314];
    assign key_original[4447] = key_shuffle[2819];
    assign key_original[4446] = key_shuffle[1512];
    assign key_original[4445] = key_shuffle[5021];
    assign key_original[4444] = key_shuffle[34];
    assign key_original[4443] = key_shuffle[4299];
    assign key_original[4442] = key_shuffle[5322];
    assign key_original[4441] = key_shuffle[3839];
    assign key_original[4440] = key_shuffle[3120];
    assign key_original[4439] = key_shuffle[4362];
    assign key_original[4438] = key_shuffle[2377];
    assign key_original[4437] = key_shuffle[1653];
    assign key_original[4436] = key_shuffle[3936];
    assign key_original[4435] = key_shuffle[544];
    assign key_original[4434] = key_shuffle[3213];
    assign key_original[4433] = key_shuffle[1216];
    assign key_original[4432] = key_shuffle[4605];
    assign key_original[4431] = key_shuffle[2915];
    assign key_original[4430] = key_shuffle[716];
    assign key_original[4429] = key_shuffle[5524];
    assign key_original[4428] = key_shuffle[4264];
    assign key_original[4427] = key_shuffle[1098];
    assign key_original[4426] = key_shuffle[2256];
    assign key_original[4425] = key_shuffle[6803];
    assign key_original[4424] = key_shuffle[3449];
    assign key_original[4423] = key_shuffle[3382];
    assign key_original[4422] = key_shuffle[404];
    assign key_original[4421] = key_shuffle[6941];
    assign key_original[4420] = key_shuffle[5456];
    assign key_original[4419] = key_shuffle[7191];
    assign key_original[4418] = key_shuffle[3698];
    assign key_original[4417] = key_shuffle[7015];
    assign key_original[4416] = key_shuffle[8095];
    assign key_original[4415] = key_shuffle[518];
    assign key_original[4414] = key_shuffle[1660];
    assign key_original[4413] = key_shuffle[4451];
    assign key_original[4412] = key_shuffle[6523];
    assign key_original[4411] = key_shuffle[6935];
    assign key_original[4410] = key_shuffle[5771];
    assign key_original[4409] = key_shuffle[1873];
    assign key_original[4408] = key_shuffle[7023];
    assign key_original[4407] = key_shuffle[319];
    assign key_original[4406] = key_shuffle[3208];
    assign key_original[4405] = key_shuffle[1754];
    assign key_original[4404] = key_shuffle[4163];
    assign key_original[4403] = key_shuffle[1289];
    assign key_original[4402] = key_shuffle[5853];
    assign key_original[4401] = key_shuffle[3409];
    assign key_original[4400] = key_shuffle[4075];
    assign key_original[4399] = key_shuffle[7216];
    assign key_original[4398] = key_shuffle[6423];
    assign key_original[4397] = key_shuffle[6869];
    assign key_original[4396] = key_shuffle[2851];
    assign key_original[4395] = key_shuffle[5130];
    assign key_original[4394] = key_shuffle[4125];
    assign key_original[4393] = key_shuffle[6243];
    assign key_original[4392] = key_shuffle[5962];
    assign key_original[4391] = key_shuffle[7171];
    assign key_original[4390] = key_shuffle[1041];
    assign key_original[4389] = key_shuffle[1833];
    assign key_original[4388] = key_shuffle[2564];
    assign key_original[4387] = key_shuffle[3699];
    assign key_original[4386] = key_shuffle[4561];
    assign key_original[4385] = key_shuffle[5936];
    assign key_original[4384] = key_shuffle[1257];
    assign key_original[4383] = key_shuffle[3758];
    assign key_original[4382] = key_shuffle[4494];
    assign key_original[4381] = key_shuffle[7615];
    assign key_original[4380] = key_shuffle[894];
    assign key_original[4379] = key_shuffle[463];
    assign key_original[4378] = key_shuffle[2711];
    assign key_original[4377] = key_shuffle[933];
    assign key_original[4376] = key_shuffle[4973];
    assign key_original[4375] = key_shuffle[2932];
    assign key_original[4374] = key_shuffle[4014];
    assign key_original[4373] = key_shuffle[192];
    assign key_original[4372] = key_shuffle[1099];
    assign key_original[4371] = key_shuffle[4020];
    assign key_original[4370] = key_shuffle[5477];
    assign key_original[4369] = key_shuffle[6106];
    assign key_original[4368] = key_shuffle[126];
    assign key_original[4367] = key_shuffle[6147];
    assign key_original[4366] = key_shuffle[7822];
    assign key_original[4365] = key_shuffle[5466];
    assign key_original[4364] = key_shuffle[6018];
    assign key_original[4363] = key_shuffle[5775];
    assign key_original[4362] = key_shuffle[3405];
    assign key_original[4361] = key_shuffle[2372];
    assign key_original[4360] = key_shuffle[2045];
    assign key_original[4359] = key_shuffle[4485];
    assign key_original[4358] = key_shuffle[5479];
    assign key_original[4357] = key_shuffle[350];
    assign key_original[4356] = key_shuffle[6555];
    assign key_original[4355] = key_shuffle[3956];
    assign key_original[4354] = key_shuffle[1078];
    assign key_original[4353] = key_shuffle[7990];
    assign key_original[4352] = key_shuffle[3436];
    assign key_original[4351] = key_shuffle[2014];
    assign key_original[4350] = key_shuffle[3743];
    assign key_original[4349] = key_shuffle[4665];
    assign key_original[4348] = key_shuffle[739];
    assign key_original[4347] = key_shuffle[233];
    assign key_original[4346] = key_shuffle[1426];
    assign key_original[4345] = key_shuffle[8190];
    assign key_original[4344] = key_shuffle[4632];
    assign key_original[4343] = key_shuffle[6693];
    assign key_original[4342] = key_shuffle[5947];
    assign key_original[4341] = key_shuffle[938];
    assign key_original[4340] = key_shuffle[2121];
    assign key_original[4339] = key_shuffle[2313];
    assign key_original[4338] = key_shuffle[8039];
    assign key_original[4337] = key_shuffle[7056];
    assign key_original[4336] = key_shuffle[3894];
    assign key_original[4335] = key_shuffle[3387];
    assign key_original[4334] = key_shuffle[1971];
    assign key_original[4333] = key_shuffle[6298];
    assign key_original[4332] = key_shuffle[8030];
    assign key_original[4331] = key_shuffle[7783];
    assign key_original[4330] = key_shuffle[4695];
    assign key_original[4329] = key_shuffle[5171];
    assign key_original[4328] = key_shuffle[6293];
    assign key_original[4327] = key_shuffle[3818];
    assign key_original[4326] = key_shuffle[5585];
    assign key_original[4325] = key_shuffle[7993];
    assign key_original[4324] = key_shuffle[7476];
    assign key_original[4323] = key_shuffle[5310];
    assign key_original[4322] = key_shuffle[4026];
    assign key_original[4321] = key_shuffle[5520];
    assign key_original[4320] = key_shuffle[3914];
    assign key_original[4319] = key_shuffle[3413];
    assign key_original[4318] = key_shuffle[1634];
    assign key_original[4317] = key_shuffle[259];
    assign key_original[4316] = key_shuffle[245];
    assign key_original[4315] = key_shuffle[744];
    assign key_original[4314] = key_shuffle[412];
    assign key_original[4313] = key_shuffle[5915];
    assign key_original[4312] = key_shuffle[3886];
    assign key_original[4311] = key_shuffle[5257];
    assign key_original[4310] = key_shuffle[7430];
    assign key_original[4309] = key_shuffle[5226];
    assign key_original[4308] = key_shuffle[3289];
    assign key_original[4307] = key_shuffle[4309];
    assign key_original[4306] = key_shuffle[7676];
    assign key_original[4305] = key_shuffle[4173];
    assign key_original[4304] = key_shuffle[5694];
    assign key_original[4303] = key_shuffle[7887];
    assign key_original[4302] = key_shuffle[1552];
    assign key_original[4301] = key_shuffle[3420];
    assign key_original[4300] = key_shuffle[6862];
    assign key_original[4299] = key_shuffle[5485];
    assign key_original[4298] = key_shuffle[4470];
    assign key_original[4297] = key_shuffle[4790];
    assign key_original[4296] = key_shuffle[4814];
    assign key_original[4295] = key_shuffle[1790];
    assign key_original[4294] = key_shuffle[4105];
    assign key_original[4293] = key_shuffle[5566];
    assign key_original[4292] = key_shuffle[5697];
    assign key_original[4291] = key_shuffle[1019];
    assign key_original[4290] = key_shuffle[5302];
    assign key_original[4289] = key_shuffle[6211];
    assign key_original[4288] = key_shuffle[2096];
    assign key_original[4287] = key_shuffle[6451];
    assign key_original[4286] = key_shuffle[3597];
    assign key_original[4285] = key_shuffle[3336];
    assign key_original[4284] = key_shuffle[7787];
    assign key_original[4283] = key_shuffle[5134];
    assign key_original[4282] = key_shuffle[1080];
    assign key_original[4281] = key_shuffle[7697];
    assign key_original[4280] = key_shuffle[763];
    assign key_original[4279] = key_shuffle[1527];
    assign key_original[4278] = key_shuffle[1151];
    assign key_original[4277] = key_shuffle[7225];
    assign key_original[4276] = key_shuffle[7229];
    assign key_original[4275] = key_shuffle[4574];
    assign key_original[4274] = key_shuffle[5780];
    assign key_original[4273] = key_shuffle[6335];
    assign key_original[4272] = key_shuffle[392];
    assign key_original[4271] = key_shuffle[4048];
    assign key_original[4270] = key_shuffle[2581];
    assign key_original[4269] = key_shuffle[7689];
    assign key_original[4268] = key_shuffle[3664];
    assign key_original[4267] = key_shuffle[2302];
    assign key_original[4266] = key_shuffle[6286];
    assign key_original[4265] = key_shuffle[6469];
    assign key_original[4264] = key_shuffle[8112];
    assign key_original[4263] = key_shuffle[3592];
    assign key_original[4262] = key_shuffle[5610];
    assign key_original[4261] = key_shuffle[6732];
    assign key_original[4260] = key_shuffle[1547];
    assign key_original[4259] = key_shuffle[3326];
    assign key_original[4258] = key_shuffle[2999];
    assign key_original[4257] = key_shuffle[7345];
    assign key_original[4256] = key_shuffle[1273];
    assign key_original[4255] = key_shuffle[4212];
    assign key_original[4254] = key_shuffle[1054];
    assign key_original[4253] = key_shuffle[5920];
    assign key_original[4252] = key_shuffle[1671];
    assign key_original[4251] = key_shuffle[7050];
    assign key_original[4250] = key_shuffle[5369];
    assign key_original[4249] = key_shuffle[4118];
    assign key_original[4248] = key_shuffle[22];
    assign key_original[4247] = key_shuffle[1205];
    assign key_original[4246] = key_shuffle[4684];
    assign key_original[4245] = key_shuffle[554];
    assign key_original[4244] = key_shuffle[3876];
    assign key_original[4243] = key_shuffle[3054];
    assign key_original[4242] = key_shuffle[5813];
    assign key_original[4241] = key_shuffle[5948];
    assign key_original[4240] = key_shuffle[7428];
    assign key_original[4239] = key_shuffle[3300];
    assign key_original[4238] = key_shuffle[5417];
    assign key_original[4237] = key_shuffle[5351];
    assign key_original[4236] = key_shuffle[1703];
    assign key_original[4235] = key_shuffle[814];
    assign key_original[4234] = key_shuffle[4630];
    assign key_original[4233] = key_shuffle[1100];
    assign key_original[4232] = key_shuffle[1275];
    assign key_original[4231] = key_shuffle[6697];
    assign key_original[4230] = key_shuffle[1601];
    assign key_original[4229] = key_shuffle[2192];
    assign key_original[4228] = key_shuffle[5288];
    assign key_original[4227] = key_shuffle[3141];
    assign key_original[4226] = key_shuffle[2137];
    assign key_original[4225] = key_shuffle[981];
    assign key_original[4224] = key_shuffle[7246];
    assign key_original[4223] = key_shuffle[444];
    assign key_original[4222] = key_shuffle[5225];
    assign key_original[4221] = key_shuffle[4628];
    assign key_original[4220] = key_shuffle[3404];
    assign key_original[4219] = key_shuffle[2699];
    assign key_original[4218] = key_shuffle[3343];
    assign key_original[4217] = key_shuffle[1370];
    assign key_original[4216] = key_shuffle[691];
    assign key_original[4215] = key_shuffle[4108];
    assign key_original[4214] = key_shuffle[502];
    assign key_original[4213] = key_shuffle[3297];
    assign key_original[4212] = key_shuffle[6476];
    assign key_original[4211] = key_shuffle[7905];
    assign key_original[4210] = key_shuffle[97];
    assign key_original[4209] = key_shuffle[7198];
    assign key_original[4208] = key_shuffle[5008];
    assign key_original[4207] = key_shuffle[848];
    assign key_original[4206] = key_shuffle[6104];
    assign key_original[4205] = key_shuffle[1398];
    assign key_original[4204] = key_shuffle[4672];
    assign key_original[4203] = key_shuffle[7470];
    assign key_original[4202] = key_shuffle[798];
    assign key_original[4201] = key_shuffle[1003];
    assign key_original[4200] = key_shuffle[6904];
    assign key_original[4199] = key_shuffle[7381];
    assign key_original[4198] = key_shuffle[6318];
    assign key_original[4197] = key_shuffle[4600];
    assign key_original[4196] = key_shuffle[386];
    assign key_original[4195] = key_shuffle[4848];
    assign key_original[4194] = key_shuffle[1780];
    assign key_original[4193] = key_shuffle[2392];
    assign key_original[4192] = key_shuffle[4987];
    assign key_original[4191] = key_shuffle[4914];
    assign key_original[4190] = key_shuffle[6402];
    assign key_original[4189] = key_shuffle[4981];
    assign key_original[4188] = key_shuffle[8163];
    assign key_original[4187] = key_shuffle[6270];
    assign key_original[4186] = key_shuffle[7163];
    assign key_original[4185] = key_shuffle[6508];
    assign key_original[4184] = key_shuffle[7442];
    assign key_original[4183] = key_shuffle[8118];
    assign key_original[4182] = key_shuffle[4421];
    assign key_original[4181] = key_shuffle[5804];
    assign key_original[4180] = key_shuffle[7071];
    assign key_original[4179] = key_shuffle[6047];
    assign key_original[4178] = key_shuffle[2743];
    assign key_original[4177] = key_shuffle[3930];
    assign key_original[4176] = key_shuffle[8108];
    assign key_original[4175] = key_shuffle[6953];
    assign key_original[4174] = key_shuffle[2402];
    assign key_original[4173] = key_shuffle[3714];
    assign key_original[4172] = key_shuffle[3852];
    assign key_original[4171] = key_shuffle[5723];
    assign key_original[4170] = key_shuffle[4878];
    assign key_original[4169] = key_shuffle[4983];
    assign key_original[4168] = key_shuffle[3489];
    assign key_original[4167] = key_shuffle[4202];
    assign key_original[4166] = key_shuffle[5309];
    assign key_original[4165] = key_shuffle[4308];
    assign key_original[4164] = key_shuffle[4527];
    assign key_original[4163] = key_shuffle[2652];
    assign key_original[4162] = key_shuffle[6900];
    assign key_original[4161] = key_shuffle[420];
    assign key_original[4160] = key_shuffle[6929];
    assign key_original[4159] = key_shuffle[3669];
    assign key_original[4158] = key_shuffle[935];
    assign key_original[4157] = key_shuffle[3659];
    assign key_original[4156] = key_shuffle[1733];
    assign key_original[4155] = key_shuffle[6348];
    assign key_original[4154] = key_shuffle[4746];
    assign key_original[4153] = key_shuffle[2515];
    assign key_original[4152] = key_shuffle[5598];
    assign key_original[4151] = key_shuffle[3801];
    assign key_original[4150] = key_shuffle[2234];
    assign key_original[4149] = key_shuffle[7083];
    assign key_original[4148] = key_shuffle[4487];
    assign key_original[4147] = key_shuffle[3983];
    assign key_original[4146] = key_shuffle[4679];
    assign key_original[4145] = key_shuffle[7607];
    assign key_original[4144] = key_shuffle[6036];
    assign key_original[4143] = key_shuffle[5794];
    assign key_original[4142] = key_shuffle[6673];
    assign key_original[4141] = key_shuffle[7480];
    assign key_original[4140] = key_shuffle[5504];
    assign key_original[4139] = key_shuffle[6281];
    assign key_original[4138] = key_shuffle[7070];
    assign key_original[4137] = key_shuffle[2481];
    assign key_original[4136] = key_shuffle[7274];
    assign key_original[4135] = key_shuffle[4279];
    assign key_original[4134] = key_shuffle[8171];
    assign key_original[4133] = key_shuffle[8147];
    assign key_original[4132] = key_shuffle[1988];
    assign key_original[4131] = key_shuffle[6180];
    assign key_original[4130] = key_shuffle[4744];
    assign key_original[4129] = key_shuffle[182];
    assign key_original[4128] = key_shuffle[7538];
    assign key_original[4127] = key_shuffle[669];
    assign key_original[4126] = key_shuffle[1832];
    assign key_original[4125] = key_shuffle[5006];
    assign key_original[4124] = key_shuffle[5442];
    assign key_original[4123] = key_shuffle[5501];
    assign key_original[4122] = key_shuffle[7157];
    assign key_original[4121] = key_shuffle[4382];
    assign key_original[4120] = key_shuffle[3968];
    assign key_original[4119] = key_shuffle[4037];
    assign key_original[4118] = key_shuffle[1088];
    assign key_original[4117] = key_shuffle[5091];
    assign key_original[4116] = key_shuffle[5755];
    assign key_original[4115] = key_shuffle[5179];
    assign key_original[4114] = key_shuffle[6500];
    assign key_original[4113] = key_shuffle[6645];
    assign key_original[4112] = key_shuffle[748];
    assign key_original[4111] = key_shuffle[1133];
    assign key_original[4110] = key_shuffle[4418];
    assign key_original[4109] = key_shuffle[6];
    assign key_original[4108] = key_shuffle[7140];
    assign key_original[4107] = key_shuffle[448];
    assign key_original[4106] = key_shuffle[6837];
    assign key_original[4105] = key_shuffle[1299];
    assign key_original[4104] = key_shuffle[4620];
    assign key_original[4103] = key_shuffle[2387];
    assign key_original[4102] = key_shuffle[4663];
    assign key_original[4101] = key_shuffle[3972];
    assign key_original[4100] = key_shuffle[7267];
    assign key_original[4099] = key_shuffle[1399];
    assign key_original[4098] = key_shuffle[7969];
    assign key_original[4097] = key_shuffle[2025];
    assign key_original[4096] = key_shuffle[2658];
    assign key_original[4095] = key_shuffle[7713];
    assign key_original[4094] = key_shuffle[4092];
    assign key_original[4093] = key_shuffle[7270];
    assign key_original[4092] = key_shuffle[5839];
    assign key_original[4091] = key_shuffle[3085];
    assign key_original[4090] = key_shuffle[1097];
    assign key_original[4089] = key_shuffle[5203];
    assign key_original[4088] = key_shuffle[7764];
    assign key_original[4087] = key_shuffle[5019];
    assign key_original[4086] = key_shuffle[1480];
    assign key_original[4085] = key_shuffle[3678];
    assign key_original[4084] = key_shuffle[2097];
    assign key_original[4083] = key_shuffle[7477];
    assign key_original[4082] = key_shuffle[8120];
    assign key_original[4081] = key_shuffle[7912];
    assign key_original[4080] = key_shuffle[4032];
    assign key_original[4079] = key_shuffle[331];
    assign key_original[4078] = key_shuffle[4888];
    assign key_original[4077] = key_shuffle[6074];
    assign key_original[4076] = key_shuffle[6340];
    assign key_original[4075] = key_shuffle[3051];
    assign key_original[4074] = key_shuffle[942];
    assign key_original[4073] = key_shuffle[585];
    assign key_original[4072] = key_shuffle[2477];
    assign key_original[4071] = key_shuffle[1979];
    assign key_original[4070] = key_shuffle[1954];
    assign key_original[4069] = key_shuffle[8003];
    assign key_original[4068] = key_shuffle[2647];
    assign key_original[4067] = key_shuffle[1340];
    assign key_original[4066] = key_shuffle[7678];
    assign key_original[4065] = key_shuffle[3766];
    assign key_original[4064] = key_shuffle[7618];
    assign key_original[4063] = key_shuffle[5313];
    assign key_original[4062] = key_shuffle[123];
    assign key_original[4061] = key_shuffle[3445];
    assign key_original[4060] = key_shuffle[220];
    assign key_original[4059] = key_shuffle[6455];
    assign key_original[4058] = key_shuffle[5418];
    assign key_original[4057] = key_shuffle[6798];
    assign key_original[4056] = key_shuffle[5998];
    assign key_original[4055] = key_shuffle[7280];
    assign key_original[4054] = key_shuffle[751];
    assign key_original[4053] = key_shuffle[5877];
    assign key_original[4052] = key_shuffle[5035];
    assign key_original[4051] = key_shuffle[2340];
    assign key_original[4050] = key_shuffle[859];
    assign key_original[4049] = key_shuffle[4664];
    assign key_original[4048] = key_shuffle[795];
    assign key_original[4047] = key_shuffle[3822];
    assign key_original[4046] = key_shuffle[3824];
    assign key_original[4045] = key_shuffle[8188];
    assign key_original[4044] = key_shuffle[7857];
    assign key_original[4043] = key_shuffle[4607];
    assign key_original[4042] = key_shuffle[2224];
    assign key_original[4041] = key_shuffle[2951];
    assign key_original[4040] = key_shuffle[438];
    assign key_original[4039] = key_shuffle[8002];
    assign key_original[4038] = key_shuffle[1406];
    assign key_original[4037] = key_shuffle[6202];
    assign key_original[4036] = key_shuffle[7459];
    assign key_original[4035] = key_shuffle[1191];
    assign key_original[4034] = key_shuffle[1266];
    assign key_original[4033] = key_shuffle[2522];
    assign key_original[4032] = key_shuffle[439];
    assign key_original[4031] = key_shuffle[3309];
    assign key_original[4030] = key_shuffle[1863];
    assign key_original[4029] = key_shuffle[2151];
    assign key_original[4028] = key_shuffle[916];
    assign key_original[4027] = key_shuffle[4879];
    assign key_original[4026] = key_shuffle[6118];
    assign key_original[4025] = key_shuffle[1184];
    assign key_original[4024] = key_shuffle[1929];
    assign key_original[4023] = key_shuffle[4969];
    assign key_original[4022] = key_shuffle[4501];
    assign key_original[4021] = key_shuffle[3851];
    assign key_original[4020] = key_shuffle[500];
    assign key_original[4019] = key_shuffle[2267];
    assign key_original[4018] = key_shuffle[4091];
    assign key_original[4017] = key_shuffle[1342];
    assign key_original[4016] = key_shuffle[7996];
    assign key_original[4015] = key_shuffle[5680];
    assign key_original[4014] = key_shuffle[2667];
    assign key_original[4013] = key_shuffle[861];
    assign key_original[4012] = key_shuffle[939];
    assign key_original[4011] = key_shuffle[3229];
    assign key_original[4010] = key_shuffle[29];
    assign key_original[4009] = key_shuffle[7800];
    assign key_original[4008] = key_shuffle[7999];
    assign key_original[4007] = key_shuffle[1462];
    assign key_original[4006] = key_shuffle[7893];
    assign key_original[4005] = key_shuffle[3979];
    assign key_original[4004] = key_shuffle[4726];
    assign key_original[4003] = key_shuffle[6971];
    assign key_original[4002] = key_shuffle[5974];
    assign key_original[4001] = key_shuffle[4232];
    assign key_original[4000] = key_shuffle[3375];
    assign key_original[3999] = key_shuffle[8173];
    assign key_original[3998] = key_shuffle[4174];
    assign key_original[3997] = key_shuffle[2351];
    assign key_original[3996] = key_shuffle[3977];
    assign key_original[3995] = key_shuffle[3159];
    assign key_original[3994] = key_shuffle[4762];
    assign key_original[3993] = key_shuffle[156];
    assign key_original[3992] = key_shuffle[3406];
    assign key_original[3991] = key_shuffle[622];
    assign key_original[3990] = key_shuffle[7991];
    assign key_original[3989] = key_shuffle[7154];
    assign key_original[3988] = key_shuffle[4711];
    assign key_original[3987] = key_shuffle[5953];
    assign key_original[3986] = key_shuffle[5370];
    assign key_original[3985] = key_shuffle[5415];
    assign key_original[3984] = key_shuffle[7126];
    assign key_original[3983] = key_shuffle[8143];
    assign key_original[3982] = key_shuffle[4142];
    assign key_original[3981] = key_shuffle[1346];
    assign key_original[3980] = key_shuffle[7959];
    assign key_original[3979] = key_shuffle[4732];
    assign key_original[3978] = key_shuffle[6163];
    assign key_original[3977] = key_shuffle[7063];
    assign key_original[3976] = key_shuffle[7333];
    assign key_original[3975] = key_shuffle[6343];
    assign key_original[3974] = key_shuffle[4330];
    assign key_original[3973] = key_shuffle[7309];
    assign key_original[3972] = key_shuffle[1761];
    assign key_original[3971] = key_shuffle[3274];
    assign key_original[3970] = key_shuffle[2378];
    assign key_original[3969] = key_shuffle[2750];
    assign key_original[3968] = key_shuffle[8092];
    assign key_original[3967] = key_shuffle[5612];
    assign key_original[3966] = key_shuffle[1104];
    assign key_original[3965] = key_shuffle[1378];
    assign key_original[3964] = key_shuffle[6380];
    assign key_original[3963] = key_shuffle[2459];
    assign key_original[3962] = key_shuffle[3986];
    assign key_original[3961] = key_shuffle[2687];
    assign key_original[3960] = key_shuffle[5076];
    assign key_original[3959] = key_shuffle[4304];
    assign key_original[3958] = key_shuffle[7539];
    assign key_original[3957] = key_shuffle[2876];
    assign key_original[3956] = key_shuffle[6782];
    assign key_original[3955] = key_shuffle[5071];
    assign key_original[3954] = key_shuffle[952];
    assign key_original[3953] = key_shuffle[2635];
    assign key_original[3952] = key_shuffle[4579];
    assign key_original[3951] = key_shuffle[6683];
    assign key_original[3950] = key_shuffle[2916];
    assign key_original[3949] = key_shuffle[3945];
    assign key_original[3948] = key_shuffle[4117];
    assign key_original[3947] = key_shuffle[5029];
    assign key_original[3946] = key_shuffle[1294];
    assign key_original[3945] = key_shuffle[5628];
    assign key_original[3944] = key_shuffle[3600];
    assign key_original[3943] = key_shuffle[7195];
    assign key_original[3942] = key_shuffle[2373];
    assign key_original[3941] = key_shuffle[2100];
    assign key_original[3940] = key_shuffle[151];
    assign key_original[3939] = key_shuffle[7031];
    assign key_original[3938] = key_shuffle[4998];
    assign key_original[3937] = key_shuffle[4241];
    assign key_original[3936] = key_shuffle[3727];
    assign key_original[3935] = key_shuffle[5108];
    assign key_original[3934] = key_shuffle[6749];
    assign key_original[3933] = key_shuffle[3464];
    assign key_original[3932] = key_shuffle[6644];
    assign key_original[3931] = key_shuffle[4352];
    assign key_original[3930] = key_shuffle[4488];
    assign key_original[3929] = key_shuffle[3570];
    assign key_original[3928] = key_shuffle[1002];
    assign key_original[3927] = key_shuffle[1831];
    assign key_original[3926] = key_shuffle[4300];
    assign key_original[3925] = key_shuffle[3860];
    assign key_original[3924] = key_shuffle[6333];
    assign key_original[3923] = key_shuffle[6685];
    assign key_original[3922] = key_shuffle[1936];
    assign key_original[3921] = key_shuffle[2305];
    assign key_original[3920] = key_shuffle[7552];
    assign key_original[3919] = key_shuffle[5162];
    assign key_original[3918] = key_shuffle[1985];
    assign key_original[3917] = key_shuffle[3014];
    assign key_original[3916] = key_shuffle[1450];
    assign key_original[3915] = key_shuffle[5890];
    assign key_original[3914] = key_shuffle[4303];
    assign key_original[3913] = key_shuffle[6169];
    assign key_original[3912] = key_shuffle[4539];
    assign key_original[3911] = key_shuffle[8059];
    assign key_original[3910] = key_shuffle[3812];
    assign key_original[3909] = key_shuffle[204];
    assign key_original[3908] = key_shuffle[1739];
    assign key_original[3907] = key_shuffle[3591];
    assign key_original[3906] = key_shuffle[4385];
    assign key_original[3905] = key_shuffle[2574];
    assign key_original[3904] = key_shuffle[6015];
    assign key_original[3903] = key_shuffle[6113];
    assign key_original[3902] = key_shuffle[1507];
    assign key_original[3901] = key_shuffle[1737];
    assign key_original[3900] = key_shuffle[5768];
    assign key_original[3899] = key_shuffle[2960];
    assign key_original[3898] = key_shuffle[6053];
    assign key_original[3897] = key_shuffle[7578];
    assign key_original[3896] = key_shuffle[3761];
    assign key_original[3895] = key_shuffle[775];
    assign key_original[3894] = key_shuffle[1940];
    assign key_original[3893] = key_shuffle[2343];
    assign key_original[3892] = key_shuffle[2985];
    assign key_original[3891] = key_shuffle[6733];
    assign key_original[3890] = key_shuffle[4877];
    assign key_original[3889] = key_shuffle[6655];
    assign key_original[3888] = key_shuffle[7250];
    assign key_original[3887] = key_shuffle[3228];
    assign key_original[3886] = key_shuffle[832];
    assign key_original[3885] = key_shuffle[1957];
    assign key_original[3884] = key_shuffle[6543];
    assign key_original[3883] = key_shuffle[7135];
    assign key_original[3882] = key_shuffle[2117];
    assign key_original[3881] = key_shuffle[3346];
    assign key_original[3880] = key_shuffle[3651];
    assign key_original[3879] = key_shuffle[5121];
    assign key_original[3878] = key_shuffle[6406];
    assign key_original[3877] = key_shuffle[3461];
    assign key_original[3876] = key_shuffle[8011];
    assign key_original[3875] = key_shuffle[2177];
    assign key_original[3874] = key_shuffle[7043];
    assign key_original[3873] = key_shuffle[1357];
    assign key_original[3872] = key_shuffle[3145];
    assign key_original[3871] = key_shuffle[1390];
    assign key_original[3870] = key_shuffle[2516];
    assign key_original[3869] = key_shuffle[7092];
    assign key_original[3868] = key_shuffle[4654];
    assign key_original[3867] = key_shuffle[4882];
    assign key_original[3866] = key_shuffle[1631];
    assign key_original[3865] = key_shuffle[285];
    assign key_original[3864] = key_shuffle[8084];
    assign key_original[3863] = key_shuffle[1497];
    assign key_original[3862] = key_shuffle[8119];
    assign key_original[3861] = key_shuffle[7320];
    assign key_original[3860] = key_shuffle[1044];
    assign key_original[3859] = key_shuffle[6069];
    assign key_original[3858] = key_shuffle[2789];
    assign key_original[3857] = key_shuffle[5910];
    assign key_original[3856] = key_shuffle[5421];
    assign key_original[3855] = key_shuffle[6133];
    assign key_original[3854] = key_shuffle[3323];
    assign key_original[3853] = key_shuffle[6044];
    assign key_original[3852] = key_shuffle[436];
    assign key_original[3851] = key_shuffle[5373];
    assign key_original[3850] = key_shuffle[475];
    assign key_original[3849] = key_shuffle[5805];
    assign key_original[3848] = key_shuffle[408];
    assign key_original[3847] = key_shuffle[6577];
    assign key_original[3846] = key_shuffle[1254];
    assign key_original[3845] = key_shuffle[8042];
    assign key_original[3844] = key_shuffle[816];
    assign key_original[3843] = key_shuffle[7200];
    assign key_original[3842] = key_shuffle[4398];
    assign key_original[3841] = key_shuffle[7708];
    assign key_original[3840] = key_shuffle[5666];
    assign key_original[3839] = key_shuffle[3116];
    assign key_original[3838] = key_shuffle[4348];
    assign key_original[3837] = key_shuffle[7845];
    assign key_original[3836] = key_shuffle[5850];
    assign key_original[3835] = key_shuffle[160];
    assign key_original[3834] = key_shuffle[1637];
    assign key_original[3833] = key_shuffle[2084];
    assign key_original[3832] = key_shuffle[4978];
    assign key_original[3831] = key_shuffle[714];
    assign key_original[3830] = key_shuffle[4096];
    assign key_original[3829] = key_shuffle[3580];
    assign key_original[3828] = key_shuffle[1312];
    assign key_original[3827] = key_shuffle[5999];
    assign key_original[3826] = key_shuffle[4731];
    assign key_original[3825] = key_shuffle[137];
    assign key_original[3824] = key_shuffle[2376];
    assign key_original[3823] = key_shuffle[808];
    assign key_original[3822] = key_shuffle[4508];
    assign key_original[3821] = key_shuffle[5040];
    assign key_original[3820] = key_shuffle[4349];
    assign key_original[3819] = key_shuffle[7716];
    assign key_original[3818] = key_shuffle[7665];
    assign key_original[3817] = key_shuffle[6627];
    assign key_original[3816] = key_shuffle[4246];
    assign key_original[3815] = key_shuffle[5219];
    assign key_original[3814] = key_shuffle[1680];
    assign key_original[3813] = key_shuffle[6338];
    assign key_original[3812] = key_shuffle[3874];
    assign key_original[3811] = key_shuffle[1146];
    assign key_original[3810] = key_shuffle[3460];
    assign key_original[3809] = key_shuffle[200];
    assign key_original[3808] = key_shuffle[4919];
    assign key_original[3807] = key_shuffle[3101];
    assign key_original[3806] = key_shuffle[1206];
    assign key_original[3805] = key_shuffle[435];
    assign key_original[3804] = key_shuffle[4823];
    assign key_original[3803] = key_shuffle[2418];
    assign key_original[3802] = key_shuffle[5333];
    assign key_original[3801] = key_shuffle[7720];
    assign key_original[3800] = key_shuffle[431];
    assign key_original[3799] = key_shuffle[7631];
    assign key_original[3798] = key_shuffle[2432];
    assign key_original[3797] = key_shuffle[2724];
    assign key_original[3796] = key_shuffle[4219];
    assign key_original[3795] = key_shuffle[5707];
    assign key_original[3794] = key_shuffle[2846];
    assign key_original[3793] = key_shuffle[209];
    assign key_original[3792] = key_shuffle[3978];
    assign key_original[3791] = key_shuffle[1016];
    assign key_original[3790] = key_shuffle[3381];
    assign key_original[3789] = key_shuffle[6671];
    assign key_original[3788] = key_shuffle[7055];
    assign key_original[3787] = key_shuffle[1366];
    assign key_original[3786] = key_shuffle[3202];
    assign key_original[3785] = key_shuffle[1106];
    assign key_original[3784] = key_shuffle[5696];
    assign key_original[3783] = key_shuffle[679];
    assign key_original[3782] = key_shuffle[6534];
    assign key_original[3781] = key_shuffle[3232];
    assign key_original[3780] = key_shuffle[4167];
    assign key_original[3779] = key_shuffle[8121];
    assign key_original[3778] = key_shuffle[4404];
    assign key_original[3777] = key_shuffle[813];
    assign key_original[3776] = key_shuffle[2018];
    assign key_original[3775] = key_shuffle[6384];
    assign key_original[3774] = key_shuffle[2174];
    assign key_original[3773] = key_shuffle[1919];
    assign key_original[3772] = key_shuffle[3451];
    assign key_original[3771] = key_shuffle[3482];
    assign key_original[3770] = key_shuffle[3707];
    assign key_original[3769] = key_shuffle[6780];
    assign key_original[3768] = key_shuffle[4234];
    assign key_original[3767] = key_shuffle[3569];
    assign key_original[3766] = key_shuffle[6696];
    assign key_original[3765] = key_shuffle[4386];
    assign key_original[3764] = key_shuffle[2891];
    assign key_original[3763] = key_shuffle[2833];
    assign key_original[3762] = key_shuffle[3729];
    assign key_original[3761] = key_shuffle[4891];
    assign key_original[3760] = key_shuffle[1109];
    assign key_original[3759] = key_shuffle[7030];
    assign key_original[3758] = key_shuffle[1819];
    assign key_original[3757] = key_shuffle[1804];
    assign key_original[3756] = key_shuffle[7372];
    assign key_original[3755] = key_shuffle[8091];
    assign key_original[3754] = key_shuffle[3567];
    assign key_original[3753] = key_shuffle[6617];
    assign key_original[3752] = key_shuffle[1520];
    assign key_original[3751] = key_shuffle[2646];
    assign key_original[3750] = key_shuffle[7307];
    assign key_original[3749] = key_shuffle[4799];
    assign key_original[3748] = key_shuffle[7601];
    assign key_original[3747] = key_shuffle[2019];
    assign key_original[3746] = key_shuffle[5807];
    assign key_original[3745] = key_shuffle[2834];
    assign key_original[3744] = key_shuffle[496];
    assign key_original[3743] = key_shuffle[7296];
    assign key_original[3742] = key_shuffle[5081];
    assign key_original[3741] = key_shuffle[4422];
    assign key_original[3740] = key_shuffle[7011];
    assign key_original[3739] = key_shuffle[2740];
    assign key_original[3738] = key_shuffle[6606];
    assign key_original[3737] = key_shuffle[5125];
    assign key_original[3736] = key_shuffle[6417];
    assign key_original[3735] = key_shuffle[6449];
    assign key_original[3734] = key_shuffle[3721];
    assign key_original[3733] = key_shuffle[2585];
    assign key_original[3732] = key_shuffle[2441];
    assign key_original[3731] = key_shuffle[6087];
    assign key_original[3730] = key_shuffle[4793];
    assign key_original[3729] = key_shuffle[6562];
    assign key_original[3728] = key_shuffle[6394];
    assign key_original[3727] = key_shuffle[3573];
    assign key_original[3726] = key_shuffle[5795];
    assign key_original[3725] = key_shuffle[4787];
    assign key_original[3724] = key_shuffle[901];
    assign key_original[3723] = key_shuffle[7484];
    assign key_original[3722] = key_shuffle[7085];
    assign key_original[3721] = key_shuffle[4468];
    assign key_original[3720] = key_shuffle[1164];
    assign key_original[3719] = key_shuffle[3426];
    assign key_original[3718] = key_shuffle[4936];
    assign key_original[3717] = key_shuffle[1229];
    assign key_original[3716] = key_shuffle[5034];
    assign key_original[3715] = key_shuffle[3339];
    assign key_original[3714] = key_shuffle[5960];
    assign key_original[3713] = key_shuffle[4302];
    assign key_original[3712] = key_shuffle[2584];
    assign key_original[3711] = key_shuffle[563];
    assign key_original[3710] = key_shuffle[1521];
    assign key_original[3709] = key_shuffle[5116];
    assign key_original[3708] = key_shuffle[5516];
    assign key_original[3707] = key_shuffle[3954];
    assign key_original[3706] = key_shuffle[711];
    assign key_original[3705] = key_shuffle[7603];
    assign key_original[3704] = key_shuffle[6212];
    assign key_original[3703] = key_shuffle[2593];
    assign key_original[3702] = key_shuffle[1813];
    assign key_original[3701] = key_shuffle[1145];
    assign key_original[3700] = key_shuffle[2230];
    assign key_original[3699] = key_shuffle[844];
    assign key_original[3698] = key_shuffle[4517];
    assign key_original[3697] = key_shuffle[4537];
    assign key_original[3696] = key_shuffle[5012];
    assign key_original[3695] = key_shuffle[7795];
    assign key_original[3694] = key_shuffle[7247];
    assign key_original[3693] = key_shuffle[2414];
    assign key_original[3692] = key_shuffle[3660];
    assign key_original[3691] = key_shuffle[3863];
    assign key_original[3690] = key_shuffle[6295];
    assign key_original[3689] = key_shuffle[6170];
    assign key_original[3688] = key_shuffle[3495];
    assign key_original[3687] = key_shuffle[4292];
    assign key_original[3686] = key_shuffle[3031];
    assign key_original[3685] = key_shuffle[4576];
    assign key_original[3684] = key_shuffle[1859];
    assign key_original[3683] = key_shuffle[7066];
    assign key_original[3682] = key_shuffle[336];
    assign key_original[3681] = key_shuffle[5816];
    assign key_original[3680] = key_shuffle[5584];
    assign key_original[3679] = key_shuffle[110];
    assign key_original[3678] = key_shuffle[3543];
    assign key_original[3677] = key_shuffle[2729];
    assign key_original[3676] = key_shuffle[4824];
    assign key_original[3675] = key_shuffle[1503];
    assign key_original[3674] = key_shuffle[3150];
    assign key_original[3673] = key_shuffle[3617];
    assign key_original[3672] = key_shuffle[2605];
    assign key_original[3671] = key_shuffle[354];
    assign key_original[3670] = key_shuffle[4283];
    assign key_original[3669] = key_shuffle[5154];
    assign key_original[3668] = key_shuffle[7730];
    assign key_original[3667] = key_shuffle[5901];
    assign key_original[3666] = key_shuffle[5186];
    assign key_original[3665] = key_shuffle[231];
    assign key_original[3664] = key_shuffle[2149];
    assign key_original[3663] = key_shuffle[4550];
    assign key_original[3662] = key_shuffle[2810];
    assign key_original[3661] = key_shuffle[5223];
    assign key_original[3660] = key_shuffle[1921];
    assign key_original[3659] = key_shuffle[1646];
    assign key_original[3658] = key_shuffle[6743];
    assign key_original[3657] = key_shuffle[6360];
    assign key_original[3656] = key_shuffle[3465];
    assign key_original[3655] = key_shuffle[4643];
    assign key_original[3654] = key_shuffle[3829];
    assign key_original[3653] = key_shuffle[2676];
    assign key_original[3652] = key_shuffle[81];
    assign key_original[3651] = key_shuffle[2175];
    assign key_original[3650] = key_shuffle[2893];
    assign key_original[3649] = key_shuffle[3612];
    assign key_original[3648] = key_shuffle[3453];
    assign key_original[3647] = key_shuffle[3648];
    assign key_original[3646] = key_shuffle[826];
    assign key_original[3645] = key_shuffle[488];
    assign key_original[3644] = key_shuffle[6596];
    assign key_original[3643] = key_shuffle[4723];
    assign key_original[3642] = key_shuffle[3384];
    assign key_original[3641] = key_shuffle[3262];
    assign key_original[3640] = key_shuffle[1086];
    assign key_original[3639] = key_shuffle[393];
    assign key_original[3638] = key_shuffle[4465];
    assign key_original[3637] = key_shuffle[5297];
    assign key_original[3636] = key_shuffle[4397];
    assign key_original[3635] = key_shuffle[5658];
    assign key_original[3634] = key_shuffle[4259];
    assign key_original[3633] = key_shuffle[4945];
    assign key_original[3632] = key_shuffle[8038];
    assign key_original[3631] = key_shuffle[7364];
    assign key_original[3630] = key_shuffle[5414];
    assign key_original[3629] = key_shuffle[4251];
    assign key_original[3628] = key_shuffle[4129];
    assign key_original[3627] = key_shuffle[3681];
    assign key_original[3626] = key_shuffle[6510];
    assign key_original[3625] = key_shuffle[5168];
    assign key_original[3624] = key_shuffle[6615];
    assign key_original[3623] = key_shuffle[4669];
    assign key_original[3622] = key_shuffle[1265];
    assign key_original[3621] = key_shuffle[4694];
    assign key_original[3620] = key_shuffle[1138];
    assign key_original[3619] = key_shuffle[7779];
    assign key_original[3618] = key_shuffle[2057];
    assign key_original[3617] = key_shuffle[3149];
    assign key_original[3616] = key_shuffle[6916];
    assign key_original[3615] = key_shuffle[3142];
    assign key_original[3614] = key_shuffle[5446];
    assign key_original[3613] = key_shuffle[5043];
    assign key_original[3612] = key_shuffle[6013];
    assign key_original[3611] = key_shuffle[5392];
    assign key_original[3610] = key_shuffle[5633];
    assign key_original[3609] = key_shuffle[2308];
    assign key_original[3608] = key_shuffle[8180];
    assign key_original[3607] = key_shuffle[6559];
    assign key_original[3606] = key_shuffle[888];
    assign key_original[3605] = key_shuffle[7134];
    assign key_original[3604] = key_shuffle[274];
    assign key_original[3603] = key_shuffle[699];
    assign key_original[3602] = key_shuffle[7728];
    assign key_original[3601] = key_shuffle[1962];
    assign key_original[3600] = key_shuffle[7776];
    assign key_original[3599] = key_shuffle[6898];
    assign key_original[3598] = key_shuffle[7850];
    assign key_original[3597] = key_shuffle[1175];
    assign key_original[3596] = key_shuffle[1102];
    assign key_original[3595] = key_shuffle[4703];
    assign key_original[3594] = key_shuffle[3795];
    assign key_original[3593] = key_shuffle[6528];
    assign key_original[3592] = key_shuffle[240];
    assign key_original[3591] = key_shuffle[1319];
    assign key_original[3590] = key_shuffle[3514];
    assign key_original[3589] = key_shuffle[6186];
    assign key_original[3588] = key_shuffle[4077];
    assign key_original[3587] = key_shuffle[7877];
    assign key_original[3586] = key_shuffle[4361];
    assign key_original[3585] = key_shuffle[1185];
    assign key_original[3584] = key_shuffle[2000];
    assign key_original[3583] = key_shuffle[6287];
    assign key_original[3582] = key_shuffle[2412];
    assign key_original[3581] = key_shuffle[2988];
    assign key_original[3580] = key_shuffle[7242];
    assign key_original[3579] = key_shuffle[289];
    assign key_original[3578] = key_shuffle[5806];
    assign key_original[3577] = key_shuffle[1898];
    assign key_original[3576] = key_shuffle[6481];
    assign key_original[3575] = key_shuffle[2503];
    assign key_original[3574] = key_shuffle[1676];
    assign key_original[3573] = key_shuffle[6458];
    assign key_original[3572] = key_shuffle[6096];
    assign key_original[3571] = key_shuffle[6130];
    assign key_original[3570] = key_shuffle[1647];
    assign key_original[3569] = key_shuffle[5060];
    assign key_original[3568] = key_shuffle[1465];
    assign key_original[3567] = key_shuffle[627];
    assign key_original[3566] = key_shuffle[7155];
    assign key_original[3565] = key_shuffle[6538];
    assign key_original[3564] = key_shuffle[6792];
    assign key_original[3563] = key_shuffle[4180];
    assign key_original[3562] = key_shuffle[575];
    assign key_original[3561] = key_shuffle[2735];
    assign key_original[3560] = key_shuffle[2610];
    assign key_original[3559] = key_shuffle[7760];
    assign key_original[3558] = key_shuffle[5852];
    assign key_original[3557] = key_shuffle[2408];
    assign key_original[3556] = key_shuffle[6713];
    assign key_original[3555] = key_shuffle[1519];
    assign key_original[3554] = key_shuffle[4315];
    assign key_original[3553] = key_shuffle[7281];
    assign key_original[3552] = key_shuffle[4031];
    assign key_original[3551] = key_shuffle[6185];
    assign key_original[3550] = key_shuffle[2770];
    assign key_original[3549] = key_shuffle[3075];
    assign key_original[3548] = key_shuffle[3329];
    assign key_original[3547] = key_shuffle[5200];
    assign key_original[3546] = key_shuffle[1415];
    assign key_original[3545] = key_shuffle[3070];
    assign key_original[3544] = key_shuffle[5595];
    assign key_original[3543] = key_shuffle[1868];
    assign key_original[3542] = key_shuffle[6504];
    assign key_original[3541] = key_shuffle[966];
    assign key_original[3540] = key_shuffle[2189];
    assign key_original[3539] = key_shuffle[5551];
    assign key_original[3538] = key_shuffle[308];
    assign key_original[3537] = key_shuffle[996];
    assign key_original[3536] = key_shuffle[3492];
    assign key_original[3535] = key_shuffle[6506];
    assign key_original[3534] = key_shuffle[293];
    assign key_original[3533] = key_shuffle[5201];
    assign key_original[3532] = key_shuffle[2452];
    assign key_original[3531] = key_shuffle[30];
    assign key_original[3530] = key_shuffle[7378];
    assign key_original[3529] = key_shuffle[2388];
    assign key_original[3528] = key_shuffle[2328];
    assign key_original[3527] = key_shuffle[4126];
    assign key_original[3526] = key_shuffle[2325];
    assign key_original[3525] = key_shuffle[5073];
    assign key_original[3524] = key_shuffle[6349];
    assign key_original[3523] = key_shuffle[4806];
    assign key_original[3522] = key_shuffle[5367];
    assign key_original[3521] = key_shuffle[7797];
    assign key_original[3520] = key_shuffle[879];
    assign key_original[3519] = key_shuffle[4638];
    assign key_original[3518] = key_shuffle[1673];
    assign key_original[3517] = key_shuffle[116];
    assign key_original[3516] = key_shuffle[717];
    assign key_original[3515] = key_shuffle[5317];
    assign key_original[3514] = key_shuffle[5590];
    assign key_original[3513] = key_shuffle[5597];
    assign key_original[3512] = key_shuffle[1705];
    assign key_original[3511] = key_shuffle[7208];
    assign key_original[3510] = key_shuffle[806];
    assign key_original[3509] = key_shuffle[6963];
    assign key_original[3508] = key_shuffle[1116];
    assign key_original[3507] = key_shuffle[3224];
    assign key_original[3506] = key_shuffle[5390];
    assign key_original[3505] = key_shuffle[1248];
    assign key_original[3504] = key_shuffle[478];
    assign key_original[3503] = key_shuffle[3443];
    assign key_original[3502] = key_shuffle[7331];
    assign key_original[3501] = key_shuffle[684];
    assign key_original[3500] = key_shuffle[372];
    assign key_original[3499] = key_shuffle[5222];
    assign key_original[3498] = key_shuffle[5957];
    assign key_original[3497] = key_shuffle[7585];
    assign key_original[3496] = key_shuffle[467];
    assign key_original[3495] = key_shuffle[3184];
    assign key_original[3494] = key_shuffle[5564];
    assign key_original[3493] = key_shuffle[2201];
    assign key_original[3492] = key_shuffle[5082];
    assign key_original[3491] = key_shuffle[2568];
    assign key_original[3490] = key_shuffle[3527];
    assign key_original[3489] = key_shuffle[6851];
    assign key_original[3488] = key_shuffle[5814];
    assign key_original[3487] = key_shuffle[6704];
    assign key_original[3486] = key_shuffle[376];
    assign key_original[3485] = key_shuffle[5228];
    assign key_original[3484] = key_shuffle[1738];
    assign key_original[3483] = key_shuffle[5996];
    assign key_original[3482] = key_shuffle[4859];
    assign key_original[3481] = key_shuffle[1559];
    assign key_original[3480] = key_shuffle[6921];
    assign key_original[3479] = key_shuffle[5410];
    assign key_original[3478] = key_shuffle[6216];
    assign key_original[3477] = key_shuffle[4984];
    assign key_original[3476] = key_shuffle[5840];
    assign key_original[3475] = key_shuffle[3506];
    assign key_original[3474] = key_shuffle[6827];
    assign key_original[3473] = key_shuffle[1327];
    assign key_original[3472] = key_shuffle[6763];
    assign key_original[3471] = key_shuffle[2031];
    assign key_original[3470] = key_shuffle[8012];
    assign key_original[3469] = key_shuffle[4556];
    assign key_original[3468] = key_shuffle[5124];
    assign key_original[3467] = key_shuffle[5172];
    assign key_original[3466] = key_shuffle[2024];
    assign key_original[3465] = key_shuffle[5329];
    assign key_original[3464] = key_shuffle[5958];
    assign key_original[3463] = key_shuffle[2494];
    assign key_original[3462] = key_shuffle[7068];
    assign key_original[3461] = key_shuffle[7878];
    assign key_original[3460] = key_shuffle[6277];
    assign key_original[3459] = key_shuffle[3062];
    assign key_original[3458] = key_shuffle[1130];
    assign key_original[3457] = key_shuffle[1746];
    assign key_original[3456] = key_shuffle[2196];
    assign key_original[3455] = key_shuffle[6363];
    assign key_original[3454] = key_shuffle[5772];
    assign key_original[3453] = key_shuffle[7666];
    assign key_original[3452] = key_shuffle[7196];
    assign key_original[3451] = key_shuffle[5026];
    assign key_original[3450] = key_shuffle[411];
    assign key_original[3449] = key_shuffle[5648];
    assign key_original[3448] = key_shuffle[7181];
    assign key_original[3447] = key_shuffle[7376];
    assign key_original[3446] = key_shuffle[2411];
    assign key_original[3445] = key_shuffle[3314];
    assign key_original[3444] = key_shuffle[6571];
    assign key_original[3443] = key_shuffle[3226];
    assign key_original[3442] = key_shuffle[4809];
    assign key_original[3441] = key_shuffle[1040];
    assign key_original[3440] = key_shuffle[1345];
    assign key_original[3439] = key_shuffle[735];
    assign key_original[3438] = key_shuffle[4042];
    assign key_original[3437] = key_shuffle[2651];
    assign key_original[3436] = key_shuffle[6404];
    assign key_original[3435] = key_shuffle[5144];
    assign key_original[3434] = key_shuffle[3825];
    assign key_original[3433] = key_shuffle[4581];
    assign key_original[3432] = key_shuffle[2198];
    assign key_original[3431] = key_shuffle[5491];
    assign key_original[3430] = key_shuffle[5603];
    assign key_original[3429] = key_shuffle[5136];
    assign key_original[3428] = key_shuffle[6059];
    assign key_original[3427] = key_shuffle[145];
    assign key_original[3426] = key_shuffle[2095];
    assign key_original[3425] = key_shuffle[5405];
    assign key_original[3424] = key_shuffle[3935];
    assign key_original[3423] = key_shuffle[6011];
    assign key_original[3422] = key_shuffle[8051];
    assign key_original[3421] = key_shuffle[5626];
    assign key_original[3420] = key_shuffle[7453];
    assign key_original[3419] = key_shuffle[1298];
    assign key_original[3418] = key_shuffle[5092];
    assign key_original[3417] = key_shuffle[6800];
    assign key_original[3416] = key_shuffle[6155];
    assign key_original[3415] = key_shuffle[4265];
    assign key_original[3414] = key_shuffle[2576];
    assign key_original[3413] = key_shuffle[1530];
    assign key_original[3412] = key_shuffle[1329];
    assign key_original[3411] = key_shuffle[5667];
    assign key_original[3410] = key_shuffle[6983];
    assign key_original[3409] = key_shuffle[4794];
    assign key_original[3408] = key_shuffle[5488];
    assign key_original[3407] = key_shuffle[5239];
    assign key_original[3406] = key_shuffle[7919];
    assign key_original[3405] = key_shuffle[8080];
    assign key_original[3404] = key_shuffle[2400];
    assign key_original[3403] = key_shuffle[6438];
    assign key_original[3402] = key_shuffle[2616];
    assign key_original[3401] = key_shuffle[4274];
    assign key_original[3400] = key_shuffle[4052];
    assign key_original[3399] = key_shuffle[682];
    assign key_original[3398] = key_shuffle[2284];
    assign key_original[3397] = key_shuffle[4082];
    assign key_original[3396] = key_shuffle[109];
    assign key_original[3395] = key_shuffle[7240];
    assign key_original[3394] = key_shuffle[5497];
    assign key_original[3393] = key_shuffle[2940];
    assign key_original[3392] = key_shuffle[2933];
    assign key_original[3391] = key_shuffle[5678];
    assign key_original[3390] = key_shuffle[6254];
    assign key_original[3389] = key_shuffle[6687];
    assign key_original[3388] = key_shuffle[1377];
    assign key_original[3387] = key_shuffle[1466];
    assign key_original[3386] = key_shuffle[5937];
    assign key_original[3385] = key_shuffle[3609];
    assign key_original[3384] = key_shuffle[5185];
    assign key_original[3383] = key_shuffle[6710];
    assign key_original[3382] = key_shuffle[2822];
    assign key_original[3381] = key_shuffle[260];
    assign key_original[3380] = key_shuffle[2691];
    assign key_original[3379] = key_shuffle[4766];
    assign key_original[3378] = key_shuffle[5924];
    assign key_original[3377] = key_shuffle[1330];
    assign key_original[3376] = key_shuffle[4093];
    assign key_original[3375] = key_shuffle[2380];
    assign key_original[3374] = key_shuffle[282];
    assign key_original[3373] = key_shuffle[5145];
    assign key_original[3372] = key_shuffle[8155];
    assign key_original[3371] = key_shuffle[2369];
    assign key_original[3370] = key_shuffle[586];
    assign key_original[3369] = key_shuffle[3282];
    assign key_original[3368] = key_shuffle[1568];
    assign key_original[3367] = key_shuffle[7889];
    assign key_original[3366] = key_shuffle[7938];
    assign key_original[3365] = key_shuffle[701];
    assign key_original[3364] = key_shuffle[4954];
    assign key_original[3363] = key_shuffle[557];
    assign key_original[3362] = key_shuffle[7120];
    assign key_original[3361] = key_shuffle[4650];
    assign key_original[3360] = key_shuffle[1743];
    assign key_original[3359] = key_shuffle[1408];
    assign key_original[3358] = key_shuffle[1468];
    assign key_original[3357] = key_shuffle[1182];
    assign key_original[3356] = key_shuffle[2363];
    assign key_original[3355] = key_shuffle[5207];
    assign key_original[3354] = key_shuffle[7550];
    assign key_original[3353] = key_shuffle[3198];
    assign key_original[3352] = key_shuffle[362];
    assign key_original[3351] = key_shuffle[1168];
    assign key_original[3350] = key_shuffle[3341];
    assign key_original[3349] = key_shuffle[1437];
    assign key_original[3348] = key_shuffle[7766];
    assign key_original[3347] = key_shuffle[3964];
    assign key_original[3346] = key_shuffle[120];
    assign key_original[3345] = key_shuffle[2803];
    assign key_original[3344] = key_shuffle[28];
    assign key_original[3343] = key_shuffle[1910];
    assign key_original[3342] = key_shuffle[3316];
    assign key_original[3341] = key_shuffle[5576];
    assign key_original[3340] = key_shuffle[3505];
    assign key_original[3339] = key_shuffle[7613];
    assign key_original[3338] = key_shuffle[4946];
    assign key_original[3337] = key_shuffle[6662];
    assign key_original[3336] = key_shuffle[4751];
    assign key_original[3335] = key_shuffle[7515];
    assign key_original[3334] = key_shuffle[2867];
    assign key_original[3333] = key_shuffle[5512];
    assign key_original[3332] = key_shuffle[7644];
    assign key_original[3331] = key_shuffle[7500];
    assign key_original[3330] = key_shuffle[8098];
    assign key_original[3329] = key_shuffle[4266];
    assign key_original[3328] = key_shuffle[510];
    assign key_original[3327] = key_shuffle[3859];
    assign key_original[3326] = key_shuffle[7415];
    assign key_original[3325] = key_shuffle[4178];
    assign key_original[3324] = key_shuffle[1153];
    assign key_original[3323] = key_shuffle[2485];
    assign key_original[3322] = key_shuffle[5242];
    assign key_original[3321] = key_shuffle[4355];
    assign key_original[3320] = key_shuffle[4081];
    assign key_original[3319] = key_shuffle[6524];
    assign key_original[3318] = key_shuffle[4231];
    assign key_original[3317] = key_shuffle[6173];
    assign key_original[3316] = key_shuffle[5917];
    assign key_original[3315] = key_shuffle[1616];
    assign key_original[3314] = key_shuffle[2027];
    assign key_original[3313] = key_shuffle[3768];
    assign key_original[3312] = key_shuffle[5718];
    assign key_original[3311] = key_shuffle[7045];
    assign key_original[3310] = key_shuffle[5631];
    assign key_original[3309] = key_shuffle[979];
    assign key_original[3308] = key_shuffle[3177];
    assign key_original[3307] = key_shuffle[3647];
    assign key_original[3306] = key_shuffle[3084];
    assign key_original[3305] = key_shuffle[2780];
    assign key_original[3304] = key_shuffle[4875];
    assign key_original[3303] = key_shuffle[5965];
    assign key_original[3302] = key_shuffle[6231];
    assign key_original[3301] = key_shuffle[567];
    assign key_original[3300] = key_shuffle[750];
    assign key_original[3299] = key_shuffle[7814];
    assign key_original[3298] = key_shuffle[4194];
    assign key_original[3297] = key_shuffle[1042];
    assign key_original[3296] = key_shuffle[934];
    assign key_original[3295] = key_shuffle[2604];
    assign key_original[3294] = key_shuffle[5511];
    assign key_original[3293] = key_shuffle[4086];
    assign key_original[3292] = key_shuffle[2521];
    assign key_original[3291] = key_shuffle[6705];
    assign key_original[3290] = key_shuffle[2124];
    assign key_original[3289] = key_shuffle[6496];
    assign key_original[3288] = key_shuffle[3294];
    assign key_original[3287] = key_shuffle[1902];
    assign key_original[3286] = key_shuffle[7433];
    assign key_original[3285] = key_shuffle[3269];
    assign key_original[3284] = key_shuffle[44];
    assign key_original[3283] = key_shuffle[1385];
    assign key_original[3282] = key_shuffle[3059];
    assign key_original[3281] = key_shuffle[5296];
    assign key_original[3280] = key_shuffle[3498];
    assign key_original[3279] = key_shuffle[6597];
    assign key_original[3278] = key_shuffle[158];
    assign key_original[3277] = key_shuffle[1434];
    assign key_original[3276] = key_shuffle[5118];
    assign key_original[3275] = key_shuffle[5744];
    assign key_original[3274] = key_shuffle[1870];
    assign key_original[3273] = key_shuffle[2913];
    assign key_original[3272] = key_shuffle[35];
    assign key_original[3271] = key_shuffle[992];
    assign key_original[3270] = key_shuffle[6146];
    assign key_original[3269] = key_shuffle[8182];
    assign key_original[3268] = key_shuffle[5070];
    assign key_original[3267] = key_shuffle[7508];
    assign key_original[3266] = key_shuffle[7105];
    assign key_original[3265] = key_shuffle[7775];
    assign key_original[3264] = key_shuffle[5261];
    assign key_original[3263] = key_shuffle[7722];
    assign key_original[3262] = key_shuffle[217];
    assign key_original[3261] = key_shuffle[8169];
    assign key_original[3260] = key_shuffle[3284];
    assign key_original[3259] = key_shuffle[1698];
    assign key_original[3258] = key_shuffle[5863];
    assign key_original[3257] = key_shuffle[6830];
    assign key_original[3256] = key_shuffle[3132];
    assign key_original[3255] = key_shuffle[1402];
    assign key_original[3254] = key_shuffle[3750];
    assign key_original[3253] = key_shuffle[3408];
    assign key_original[3252] = key_shuffle[3480];
    assign key_original[3251] = key_shuffle[7373];
    assign key_original[3250] = key_shuffle[1347];
    assign key_original[3249] = key_shuffle[4874];
    assign key_original[3248] = key_shuffle[1306];
    assign key_original[3247] = key_shuffle[2475];
    assign key_original[3246] = key_shuffle[6296];
    assign key_original[3245] = key_shuffle[1759];
    assign key_original[3244] = key_shuffle[4275];
    assign key_original[3243] = key_shuffle[6150];
    assign key_original[3242] = key_shuffle[4640];
    assign key_original[3241] = key_shuffle[2422];
    assign key_original[3240] = key_shuffle[647];
    assign key_original[3239] = key_shuffle[6518];
    assign key_original[3238] = key_shuffle[1794];
    assign key_original[3237] = key_shuffle[3985];
    assign key_original[3236] = key_shuffle[1846];
    assign key_original[3235] = key_shuffle[7598];
    assign key_original[3234] = key_shuffle[348];
    assign key_original[3233] = key_shuffle[963];
    assign key_original[3232] = key_shuffle[5249];
    assign key_original[3231] = key_shuffle[1063];
    assign key_original[3230] = key_shuffle[3971];
    assign key_original[3229] = key_shuffle[1719];
    assign key_original[3228] = key_shuffle[4635];
    assign key_original[3227] = key_shuffle[2637];
    assign key_original[3226] = key_shuffle[7920];
    assign key_original[3225] = key_shuffle[1667];
    assign key_original[3224] = key_shuffle[779];
    assign key_original[3223] = key_shuffle[3807];
    assign key_original[3222] = key_shuffle[4000];
    assign key_original[3221] = key_shuffle[6919];
    assign key_original[3220] = key_shuffle[4943];
    assign key_original[3219] = key_shuffle[650];
    assign key_original[3218] = key_shuffle[6646];
    assign key_original[3217] = key_shuffle[3454];
    assign key_original[3216] = key_shuffle[2029];
    assign key_original[3215] = key_shuffle[5686];
    assign key_original[3214] = key_shuffle[6840];
    assign key_original[3213] = key_shuffle[3136];
    assign key_original[3212] = key_shuffle[5235];
    assign key_original[3211] = key_shuffle[6668];
    assign key_original[3210] = key_shuffle[6446];
    assign key_original[3209] = key_shuffle[1994];
    assign key_original[3208] = key_shuffle[5065];
    assign key_original[3207] = key_shuffle[4150];
    assign key_original[3206] = key_shuffle[3552];
    assign key_original[3205] = key_shuffle[2723];
    assign key_original[3204] = key_shuffle[4785];
    assign key_original[3203] = key_shuffle[2598];
    assign key_original[3202] = key_shuffle[7310];
    assign key_original[3201] = key_shuffle[1361];
    assign key_original[3200] = key_shuffle[5476];
    assign key_original[3199] = key_shuffle[1650];
    assign key_original[3198] = key_shuffle[6426];
    assign key_original[3197] = key_shuffle[3740];
    assign key_original[3196] = key_shuffle[3338];
    assign key_original[3195] = key_shuffle[6285];
    assign key_original[3194] = key_shuffle[7213];
    assign key_original[3193] = key_shuffle[7929];
    assign key_original[3192] = key_shuffle[818];
    assign key_original[3191] = key_shuffle[4354];
    assign key_original[3190] = key_shuffle[1028];
    assign key_original[3189] = key_shuffle[828];
    assign key_original[3188] = key_shuffle[2697];
    assign key_original[3187] = key_shuffle[3776];
    assign key_original[3186] = key_shuffle[4267];
    assign key_original[3185] = key_shuffle[7254];
    assign key_original[3184] = key_shuffle[1120];
    assign key_original[3183] = key_shuffle[5879];
    assign key_original[3182] = key_shuffle[458];
    assign key_original[3181] = key_shuffle[5664];
    assign key_original[3180] = key_shuffle[2370];
    assign key_original[3179] = key_shuffle[1325];
    assign key_original[3178] = key_shuffle[8006];
    assign key_original[3177] = key_shuffle[3433];
    assign key_original[3176] = key_shuffle[4104];
    assign key_original[3175] = key_shuffle[8018];
    assign key_original[3174] = key_shuffle[6324];
    assign key_original[3173] = key_shuffle[4384];
    assign key_original[3172] = key_shuffle[5919];
    assign key_original[3171] = key_shuffle[2898];
    assign key_original[3170] = key_shuffle[4775];
    assign key_original[3169] = key_shuffle[7393];
    assign key_original[3168] = key_shuffle[6968];
    assign key_original[3167] = key_shuffle[990];
    assign key_original[3166] = key_shuffle[2339];
    assign key_original[3165] = key_shuffle[2479];
    assign key_original[3164] = key_shuffle[3806];
    assign key_original[3163] = key_shuffle[5698];
    assign key_original[3162] = key_shuffle[5075];
    assign key_original[3161] = key_shuffle[2120];
    assign key_original[3160] = key_shuffle[15];
    assign key_original[3159] = key_shuffle[8181];
    assign key_original[3158] = key_shuffle[5928];
    assign key_original[3157] = key_shuffle[8028];
    assign key_original[3156] = key_shuffle[2532];
    assign key_original[3155] = key_shuffle[1543];
    assign key_original[3154] = key_shuffle[5018];
    assign key_original[3153] = key_shuffle[8116];
    assign key_original[3152] = key_shuffle[6591];
    assign key_original[3151] = key_shuffle[2950];
    assign key_original[3150] = key_shuffle[928];
    assign key_original[3149] = key_shuffle[5724];
    assign key_original[3148] = key_shuffle[4217];
    assign key_original[3147] = key_shuffle[2265];
    assign key_original[3146] = key_shuffle[7736];
    assign key_original[3145] = key_shuffle[3504];
    assign key_original[3144] = key_shuffle[2219];
    assign key_original[3143] = key_shuffle[3354];
    assign key_original[3142] = key_shuffle[2135];
    assign key_original[3141] = key_shuffle[671];
    assign key_original[3140] = key_shuffle[2688];
    assign key_original[3139] = key_shuffle[1630];
    assign key_original[3138] = key_shuffle[1224];
    assign key_original[3137] = key_shuffle[4957];
    assign key_original[3136] = key_shuffle[5635];
    assign key_original[3135] = key_shuffle[265];
    assign key_original[3134] = key_shuffle[6509];
    assign key_original[3133] = key_shuffle[4346];
    assign key_original[3132] = key_shuffle[3473];
    assign key_original[3131] = key_shuffle[1854];
    assign key_original[3130] = key_shuffle[4288];
    assign key_original[3129] = key_shuffle[5428];
    assign key_original[3128] = key_shuffle[5182];
    assign key_original[3127] = key_shuffle[3363];
    assign key_original[3126] = key_shuffle[2736];
    assign key_original[3125] = key_shuffle[5844];
    assign key_original[3124] = key_shuffle[1010];
    assign key_original[3123] = key_shuffle[4238];
    assign key_original[3122] = key_shuffle[3838];
    assign key_original[3121] = key_shuffle[4497];
    assign key_original[3120] = key_shuffle[55];
    assign key_original[3119] = key_shuffle[5864];
    assign key_original[3118] = key_shuffle[3187];
    assign key_original[3117] = key_shuffle[5160];
    assign key_original[3116] = key_shuffle[326];
    assign key_original[3115] = key_shuffle[1252];
    assign key_original[3114] = key_shuffle[6444];
    assign key_original[3113] = key_shuffle[286];
    assign key_original[3112] = key_shuffle[3172];
    assign key_original[3111] = key_shuffle[205];
    assign key_original[3110] = key_shuffle[6120];
    assign key_original[3109] = key_shuffle[686];
    assign key_original[3108] = key_shuffle[5212];
    assign key_original[3107] = key_shuffle[2279];
    assign key_original[3106] = key_shuffle[5854];
    assign key_original[3105] = key_shuffle[2733];
    assign key_original[3104] = key_shuffle[3677];
    assign key_original[3103] = key_shuffle[4034];
    assign key_original[3102] = key_shuffle[1196];
    assign key_original[3101] = key_shuffle[3836];
    assign key_original[3100] = key_shuffle[7568];
    assign key_original[3099] = key_shuffle[2405];
    assign key_original[3098] = key_shuffle[6051];
    assign key_original[3097] = key_shuffle[7981];
    assign key_original[3096] = key_shuffle[3458];
    assign key_original[3095] = key_shuffle[7451];
    assign key_original[3094] = key_shuffle[956];
    assign key_original[3093] = key_shuffle[5872];
    assign key_original[3092] = key_shuffle[824];
    assign key_original[3091] = key_shuffle[304];
    assign key_original[3090] = key_shuffle[5607];
    assign key_original[3089] = key_shuffle[7677];
    assign key_original[3088] = key_shuffle[2033];
    assign key_original[3087] = key_shuffle[4992];
    assign key_original[3086] = key_shuffle[2748];
    assign key_original[3085] = key_shuffle[5539];
    assign key_original[3084] = key_shuffle[5334];
    assign key_original[3083] = key_shuffle[5577];
    assign key_original[3082] = key_shuffle[8015];
    assign key_original[3081] = key_shuffle[4254];
    assign key_original[3080] = key_shuffle[2107];
    assign key_original[3079] = key_shuffle[4029];
    assign key_original[3078] = key_shuffle[719];
    assign key_original[3077] = key_shuffle[1883];
    assign key_original[3076] = key_shuffle[7695];
    assign key_original[3075] = key_shuffle[4380];
    assign key_original[3074] = key_shuffle[7016];
    assign key_original[3073] = key_shuffle[1351];
    assign key_original[3072] = key_shuffle[3666];
    assign key_original[3071] = key_shuffle[7939];
    assign key_original[3070] = key_shuffle[329];
    assign key_original[3069] = key_shuffle[1751];
    assign key_original[3068] = key_shuffle[6726];
    assign key_original[3067] = key_shuffle[2690];
    assign key_original[3066] = key_shuffle[4196];
    assign key_original[3065] = key_shuffle[7308];
    assign key_original[3064] = key_shuffle[5085];
    assign key_original[3063] = key_shuffle[5153];
    assign key_original[3062] = key_shuffle[8094];
    assign key_original[3061] = key_shuffle[2386];
    assign key_original[3060] = key_shuffle[1890];
    assign key_original[3059] = key_shuffle[7512];
    assign key_original[3058] = key_shuffle[2903];
    assign key_original[3057] = key_shuffle[6308];
    assign key_original[3056] = key_shuffle[4467];
    assign key_original[3055] = key_shuffle[7583];
    assign key_original[3054] = key_shuffle[3374];
    assign key_original[3053] = key_shuffle[3121];
    assign key_original[3052] = key_shuffle[7582];
    assign key_original[3051] = key_shuffle[3779];
    assign key_original[3050] = key_shuffle[2558];
    assign key_original[3049] = key_shuffle[4720];
    assign key_original[3048] = key_shuffle[2509];
    assign key_original[3047] = key_shuffle[6090];
    assign key_original[3046] = key_shuffle[1166];
    assign key_original[3045] = key_shuffle[2315];
    assign key_original[3044] = key_shuffle[7590];
    assign key_original[3043] = key_shuffle[6403];
    assign key_original[3042] = key_shuffle[4662];
    assign key_original[3041] = key_shuffle[4004];
    assign key_original[3040] = key_shuffle[7493];
    assign key_original[3039] = key_shuffle[4991];
    assign key_original[3038] = key_shuffle[3468];
    assign key_original[3037] = key_shuffle[2266];
    assign key_original[3036] = key_shuffle[3938];
    assign key_original[3035] = key_shuffle[4145];
    assign key_original[3034] = key_shuffle[6502];
    assign key_original[3033] = key_shuffle[1127];
    assign key_original[3032] = key_shuffle[7592];
    assign key_original[3031] = key_shuffle[1424];
    assign key_original[3030] = key_shuffle[4512];
    assign key_original[3029] = key_shuffle[4054];
    assign key_original[3028] = key_shuffle[6894];
    assign key_original[3027] = key_shuffle[8107];
    assign key_original[3026] = key_shuffle[277];
    assign key_original[3025] = key_shuffle[7562];
    assign key_original[3024] = key_shuffle[1341];
    assign key_original[3023] = key_shuffle[8065];
    assign key_original[3022] = key_shuffle[6079];
    assign key_original[3021] = key_shuffle[3035];
    assign key_original[3020] = key_shuffle[4827];
    assign key_original[3019] = key_shuffle[2104];
    assign key_original[3018] = key_shuffle[6204];
    assign key_original[3017] = key_shuffle[6187];
    assign key_original[3016] = key_shuffle[1861];
    assign key_original[3015] = key_shuffle[3809];
    assign key_original[3014] = key_shuffle[690];
    assign key_original[3013] = key_shuffle[1903];
    assign key_original[3012] = key_shuffle[3096];
    assign key_original[3011] = key_shuffle[6709];
    assign key_original[3010] = key_shuffle[7119];
    assign key_original[3009] = key_shuffle[5581];
    assign key_original[3008] = key_shuffle[850];
    assign key_original[3007] = key_shuffle[5058];
    assign key_original[3006] = key_shuffle[3053];
    assign key_original[3005] = key_shuffle[5117];
    assign key_original[3004] = key_shuffle[7125];
    assign key_original[3003] = key_shuffle[1872];
    assign key_original[3002] = key_shuffle[6873];
    assign key_original[3001] = key_shuffle[4858];
    assign key_original[3000] = key_shuffle[1004];
    assign key_original[2999] = key_shuffle[4375];
    assign key_original[2998] = key_shuffle[6356];
    assign key_original[2997] = key_shuffle[7806];
    assign key_original[2996] = key_shuffle[1343];
    assign key_original[2995] = key_shuffle[1874];
    assign key_original[2994] = key_shuffle[7837];
    assign key_original[2993] = key_shuffle[7305];
    assign key_original[2992] = key_shuffle[1588];
    assign key_original[2991] = key_shuffle[1986];
    assign key_original[2990] = key_shuffle[2957];
    assign key_original[2989] = key_shuffle[4840];
    assign key_original[2988] = key_shuffle[3371];
    assign key_original[2987] = key_shuffle[7860];
    assign key_original[2986] = key_shuffle[991];
    assign key_original[2985] = key_shuffle[5978];
    assign key_original[2984] = key_shuffle[1352];
    assign key_original[2983] = key_shuffle[4844];
    assign key_original[2982] = key_shuffle[7184];
    assign key_original[2981] = key_shuffle[3821];
    assign key_original[2980] = key_shuffle[5005];
    assign key_original[2979] = key_shuffle[5234];
    assign key_original[2978] = key_shuffle[6747];
    assign key_original[2977] = key_shuffle[7683];
    assign key_original[2976] = key_shuffle[5030];
    assign key_original[2975] = key_shuffle[2092];
    assign key_original[2974] = key_shuffle[7337];
    assign key_original[2973] = key_shuffle[4609];
    assign key_original[2972] = key_shuffle[2480];
    assign key_original[2971] = key_shuffle[2254];
    assign key_original[2970] = key_shuffle[1217];
    assign key_original[2969] = key_shuffle[6505];
    assign key_original[2968] = key_shuffle[7526];
    assign key_original[2967] = key_shuffle[7958];
    assign key_original[2966] = key_shuffle[364];
    assign key_original[2965] = key_shuffle[2620];
    assign key_original[2964] = key_shuffle[4423];
    assign key_original[2963] = key_shuffle[3638];
    assign key_original[2962] = key_shuffle[4013];
    assign key_original[2961] = key_shuffle[2941];
    assign key_original[2960] = key_shuffle[5264];
    assign key_original[2959] = key_shuffle[2471];
    assign key_original[2958] = key_shuffle[4592];
    assign key_original[2957] = key_shuffle[643];
    assign key_original[2956] = key_shuffle[7542];
    assign key_original[2955] = key_shuffle[494];
    assign key_original[2954] = key_shuffle[2732];
    assign key_original[2953] = key_shuffle[3238];
    assign key_original[2952] = key_shuffle[6138];
    assign key_original[2951] = key_shuffle[7330];
    assign key_original[2950] = key_shuffle[5907];
    assign key_original[2949] = key_shuffle[1644];
    assign key_original[2948] = key_shuffle[1684];
    assign key_original[2947] = key_shuffle[2871];
    assign key_original[2946] = key_shuffle[294];
    assign key_original[2945] = key_shuffle[2026];
    assign key_original[2944] = key_shuffle[1397];
    assign key_original[2943] = key_shuffle[234];
    assign key_original[2942] = key_shuffle[7481];
    assign key_original[2941] = key_shuffle[2887];
    assign key_original[2940] = key_shuffle[5800];
    assign key_original[2939] = key_shuffle[7434];
    assign key_original[2938] = key_shuffle[1901];
    assign key_original[2937] = key_shuffle[1964];
    assign key_original[2936] = key_shuffle[3126];
    assign key_original[2935] = key_shuffle[1457];
    assign key_original[2934] = key_shuffle[1967];
    assign key_original[2933] = key_shuffle[2683];
    assign key_original[2932] = key_shuffle[7749];
    assign key_original[2931] = key_shuffle[1034];
    assign key_original[2930] = key_shuffle[5490];
    assign key_original[2929] = key_shuffle[5208];
    assign key_original[2928] = key_shuffle[3439];
    assign key_original[2927] = key_shuffle[2506];
    assign key_original[2926] = key_shuffle[1409];
    assign key_original[2925] = key_shuffle[7807];
    assign key_original[2924] = key_shuffle[633];
    assign key_original[2923] = key_shuffle[7093];
    assign key_original[2922] = key_shuffle[6109];
    assign key_original[2921] = key_shuffle[7122];
    assign key_original[2920] = key_shuffle[75];
    assign key_original[2919] = key_shuffle[736];
    assign key_original[2918] = key_shuffle[7659];
    assign key_original[2917] = key_shuffle[4478];
    assign key_original[2916] = key_shuffle[4558];
    assign key_original[2915] = key_shuffle[1791];
    assign key_original[2914] = key_shuffle[5440];
    assign key_original[2913] = key_shuffle[6897];
    assign key_original[2912] = key_shuffle[6985];
    assign key_original[2911] = key_shuffle[3216];
    assign key_original[2910] = key_shuffle[7742];
    assign key_original[2909] = key_shuffle[4829];
    assign key_original[2908] = key_shuffle[48];
    assign key_original[2907] = key_shuffle[4440];
    assign key_original[2906] = key_shuffle[3260];
    assign key_original[2905] = key_shuffle[4866];
    assign key_original[2904] = key_shuffle[3010];
    assign key_original[2903] = key_shuffle[1679];
    assign key_original[2902] = key_shuffle[135];
    assign key_original[2901] = key_shuffle[1364];
    assign key_original[2900] = key_shuffle[7726];
    assign key_original[2899] = key_shuffle[6622];
    assign key_original[2898] = key_shuffle[4700];
    assign key_original[2897] = key_shuffle[4166];
    assign key_original[2896] = key_shuffle[4677];
    assign key_original[2895] = key_shuffle[603];
    assign key_original[2894] = key_shuffle[3913];
    assign key_original[2893] = key_shuffle[3093];
    assign key_original[2892] = key_shuffle[4963];
    assign key_original[2891] = key_shuffle[5519];
    assign key_original[2890] = key_shuffle[5695];
    assign key_original[2889] = key_shuffle[656];
    assign key_original[2888] = key_shuffle[6984];
    assign key_original[2887] = key_shuffle[5109];
    assign key_original[2886] = key_shuffle[7223];
    assign key_original[2885] = key_shuffle[5244];
    assign key_original[2884] = key_shuffle[6969];
    assign key_original[2883] = key_shuffle[1237];
    assign key_original[2882] = key_shuffle[5448];
    assign key_original[2881] = key_shuffle[357];
    assign key_original[2880] = key_shuffle[403];
    assign key_original[2879] = key_shuffle[3671];
    assign key_original[2878] = key_shuffle[6358];
    assign key_original[2877] = key_shuffle[6045];
    assign key_original[2876] = key_shuffle[6378];
    assign key_original[2875] = key_shuffle[5336];
    assign key_original[2874] = key_shuffle[2744];
    assign key_original[2873] = key_shuffle[2580];
    assign key_original[2872] = key_shuffle[2553];
    assign key_original[2871] = key_shuffle[6681];
    assign key_original[2870] = key_shuffle[944];
    assign key_original[2869] = key_shuffle[4573];
    assign key_original[2868] = key_shuffle[2542];
    assign key_original[2867] = key_shuffle[2601];
    assign key_original[2866] = key_shuffle[2694];
    assign key_original[2865] = key_shuffle[3709];
    assign key_original[2864] = key_shuffle[5973];
    assign key_original[2863] = key_shuffle[13];
    assign key_original[2862] = key_shuffle[5860];
    assign key_original[2861] = key_shuffle[7701];
    assign key_original[2860] = key_shuffle[4012];
    assign key_original[2859] = key_shuffle[430];
    assign key_original[2858] = key_shuffle[5435];
    assign key_original[2857] = key_shuffle[1848];
    assign key_original[2856] = key_shuffle[2882];
    assign key_original[2855] = key_shuffle[3013];
    assign key_original[2854] = key_shuffle[4008];
    assign key_original[2853] = key_shuffle[4323];
    assign key_original[2852] = key_shuffle[7732];
    assign key_original[2851] = key_shuffle[2706];
    assign key_original[2850] = key_shuffle[7275];
    assign key_original[2849] = key_shuffle[900];
    assign key_original[2848] = key_shuffle[7804];
    assign key_original[2847] = key_shuffle[5604];
    assign key_original[2846] = key_shuffle[7463];
    assign key_original[2845] = key_shuffle[2629];
    assign key_original[2844] = key_shuffle[46];
    assign key_original[2843] = key_shuffle[4968];
    assign key_original[2842] = key_shuffle[6989];
    assign key_original[2841] = key_shuffle[70];
    assign key_original[2840] = key_shuffle[7874];
    assign key_original[2839] = key_shuffle[6910];
    assign key_original[2838] = key_shuffle[1583];
    assign key_original[2837] = key_shuffle[8010];
    assign key_original[2836] = key_shuffle[5389];
    assign key_original[2835] = key_shuffle[3192];
    assign key_original[2834] = key_shuffle[3996];
    assign key_original[2833] = key_shuffle[7257];
    assign key_original[2832] = key_shuffle[3837];
    assign key_original[2831] = key_shuffle[3025];
    assign key_original[2830] = key_shuffle[5080];
    assign key_original[2829] = key_shuffle[2232];
    assign key_original[2828] = key_shuffle[2665];
    assign key_original[2827] = key_shuffle[187];
    assign key_original[2826] = key_shuffle[2543];
    assign key_original[2825] = key_shuffle[3526];
    assign key_original[2824] = key_shuffle[1211];
    assign key_original[2823] = key_shuffle[1015];
    assign key_original[2822] = key_shuffle[8004];
    assign key_original[2821] = key_shuffle[2345];
    assign key_original[2820] = key_shuffle[4058];
    assign key_original[2819] = key_shuffle[6354];
    assign key_original[2818] = key_shuffle[3317];
    assign key_original[2817] = key_shuffle[681];
    assign key_original[2816] = key_shuffle[5976];
    assign key_original[2815] = key_shuffle[7432];
    assign key_original[2814] = key_shuffle[6017];
    assign key_original[2813] = key_shuffle[6305];
    assign key_original[2812] = key_shuffle[3622];
    assign key_original[2811] = key_shuffle[7054];
    assign key_original[2810] = key_shuffle[7420];
    assign key_original[2809] = key_shuffle[6290];
    assign key_original[2808] = key_shuffle[5379];
    assign key_original[2807] = key_shuffle[3958];
    assign key_original[2806] = key_shuffle[1735];
    assign key_original[2805] = key_shuffle[2383];
    assign key_original[2804] = key_shuffle[2004];
    assign key_original[2803] = key_shuffle[4023];
    assign key_original[2802] = key_shuffle[2281];
    assign key_original[2801] = key_shuffle[5777];
    assign key_original[2800] = key_shuffle[1857];
    assign key_original[2799] = key_shuffle[5935];
    assign key_original[2798] = key_shuffle[6077];
    assign key_original[2797] = key_shuffle[7645];
    assign key_original[2796] = key_shuffle[7844];
    assign key_original[2795] = key_shuffle[7350];
    assign key_original[2794] = key_shuffle[3042];
    assign key_original[2793] = key_shuffle[5653];
    assign key_original[2792] = key_shuffle[3654];
    assign key_original[2791] = key_shuffle[4015];
    assign key_original[2790] = key_shuffle[1708];
    assign key_original[2789] = key_shuffle[4215];
    assign key_original[2788] = key_shuffle[4930];
    assign key_original[2787] = key_shuffle[4197];
    assign key_original[2786] = key_shuffle[6856];
    assign key_original[2785] = key_shuffle[5550];
    assign key_original[2784] = key_shuffle[2356];
    assign key_original[2783] = key_shuffle[1717];
    assign key_original[2782] = key_shuffle[1478];
    assign key_original[2781] = key_shuffle[6533];
    assign key_original[2780] = key_shuffle[437];
    assign key_original[2779] = key_shuffle[6667];
    assign key_original[2778] = key_shuffle[7017];
    assign key_original[2777] = key_shuffle[3414];
    assign key_original[2776] = key_shuffle[615];
    assign key_original[2775] = key_shuffle[2679];
    assign key_original[2774] = key_shuffle[6934];
    assign key_original[2773] = key_shuffle[1048];
    assign key_original[2772] = key_shuffle[4324];
    assign key_original[2771] = key_shuffle[5711];
    assign key_original[2770] = key_shuffle[7548];
    assign key_original[2769] = key_shuffle[36];
    assign key_original[2768] = key_shuffle[5105];
    assign key_original[2767] = key_shuffle[1563];
    assign key_original[2766] = key_shuffle[5544];
    assign key_original[2765] = key_shuffle[184];
    assign key_original[2764] = key_shuffle[7802];
    assign key_original[2763] = key_shuffle[5846];
    assign key_original[2762] = key_shuffle[4412];
    assign key_original[2761] = key_shuffle[569];
    assign key_original[2760] = key_shuffle[2264];
    assign key_original[2759] = key_shuffle[3742];
    assign key_original[2758] = key_shuffle[4314];
    assign key_original[2757] = key_shuffle[2488];
    assign key_original[2756] = key_shuffle[4952];
    assign key_original[2755] = key_shuffle[6694];
    assign key_original[2754] = key_shuffle[2258];
    assign key_original[2753] = key_shuffle[5057];
    assign key_original[2752] = key_shuffle[5123];
    assign key_original[2751] = key_shuffle[6164];
    assign key_original[2750] = key_shuffle[4755];
    assign key_original[2749] = key_shuffle[8150];
    assign key_original[2748] = key_shuffle[6352];
    assign key_original[2747] = key_shuffle[4658];
    assign key_original[2746] = key_shuffle[5184];
    assign key_original[2745] = key_shuffle[5365];
    assign key_original[2744] = key_shuffle[3683];
    assign key_original[2743] = key_shuffle[37];
    assign key_original[2742] = key_shuffle[5181];
    assign key_original[2741] = key_shuffle[4813];
    assign key_original[2740] = key_shuffle[6501];
    assign key_original[2739] = key_shuffle[5847];
    assign key_original[2738] = key_shuffle[256];
    assign key_original[2737] = key_shuffle[3325];
    assign key_original[2736] = key_shuffle[4345];
    assign key_original[2735] = key_shuffle[7757];
    assign key_original[2734] = key_shuffle[825];
    assign key_original[2733] = key_shuffle[1060];
    assign key_original[2732] = key_shuffle[7006];
    assign key_original[2731] = key_shuffle[1687];
    assign key_original[2730] = key_shuffle[758];
    assign key_original[2729] = key_shuffle[6278];
    assign key_original[2728] = key_shuffle[8072];
    assign key_original[2727] = key_shuffle[7359];
    assign key_original[2726] = key_shuffle[7355];
    assign key_original[2725] = key_shuffle[4934];
    assign key_original[2724] = key_shuffle[5246];
    assign key_original[2723] = key_shuffle[4652];
    assign key_original[2722] = key_shuffle[6607];
    assign key_original[2721] = key_shuffle[3944];
    assign key_original[2720] = key_shuffle[391];
    assign key_original[2719] = key_shuffle[5299];
    assign key_original[2718] = key_shuffle[2812];
    assign key_original[2717] = key_shuffle[6729];
    assign key_original[2716] = key_shuffle[3170];
    assign key_original[2715] = key_shuffle[803];
    assign key_original[2714] = key_shuffle[620];
    assign key_original[2713] = key_shuffle[2873];
    assign key_original[2712] = key_shuffle[2783];
    assign key_original[2711] = key_shuffle[727];
    assign key_original[2710] = key_shuffle[2767];
    assign key_original[2709] = key_shuffle[7110];
    assign key_original[2708] = key_shuffle[2978];
    assign key_original[2707] = key_shuffle[6720];
    assign key_original[2706] = key_shuffle[4405];
    assign key_original[2705] = key_shuffle[2083];
    assign key_original[2704] = key_shuffle[4956];
    assign key_original[2703] = key_shuffle[4410];
    assign key_original[2702] = key_shuffle[2429];
    assign key_original[2701] = key_shuffle[226];
    assign key_original[2700] = key_shuffle[4185];
    assign key_original[2699] = key_shuffle[8047];
    assign key_original[2698] = key_shuffle[6184];
    assign key_original[2697] = key_shuffle[5292];
    assign key_original[2696] = key_shuffle[2888];
    assign key_original[2695] = key_shuffle[2984];
    assign key_original[2694] = key_shuffle[2906];
    assign key_original[2693] = key_shuffle[1577];
    assign key_original[2692] = key_shuffle[5217];
    assign key_original[2691] = key_shuffle[2211];
    assign key_original[2690] = key_shuffle[5661];
    assign key_original[2689] = key_shuffle[4073];
    assign key_original[2688] = key_shuffle[221];
    assign key_original[2687] = key_shuffle[5922];
    assign key_original[2686] = key_shuffle[6198];
    assign key_original[2685] = key_shuffle[2011];
    assign key_original[2684] = key_shuffle[4239];
    assign key_original[2683] = key_shuffle[5783];
    assign key_original[2682] = key_shuffle[2442];
    assign key_original[2681] = key_shuffle[7144];
    assign key_original[2680] = key_shuffle[534];
    assign key_original[2679] = key_shuffle[276];
    assign key_original[2678] = key_shuffle[5355];
    assign key_original[2677] = key_shuffle[3616];
    assign key_original[2676] = key_shuffle[662];
    assign key_original[2675] = key_shuffle[7770];
    assign key_original[2674] = key_shuffle[4395];
    assign key_original[2673] = key_shuffle[5106];
    assign key_original[2672] = key_shuffle[855];
    assign key_original[2671] = key_shuffle[3834];
    assign key_original[2670] = key_shuffle[3572];
    assign key_original[2669] = key_shuffle[5174];
    assign key_original[2668] = key_shuffle[5567];
    assign key_original[2667] = key_shuffle[423];
    assign key_original[2666] = key_shuffle[1803];
    assign key_original[2665] = key_shuffle[7627];
    assign key_original[2664] = key_shuffle[7788];
    assign key_original[2663] = key_shuffle[1101];
    assign key_original[2662] = key_shuffle[2087];
    assign key_original[2661] = key_shuffle[3631];
    assign key_original[2660] = key_shuffle[347];
    assign key_original[2659] = key_shuffle[2098];
    assign key_original[2658] = key_shuffle[5732];
    assign key_original[2657] = key_shuffle[7835];
    assign key_original[2656] = key_shuffle[3895];
    assign key_original[2655] = key_shuffle[7033];
    assign key_original[2654] = key_shuffle[3474];
    assign key_original[2653] = key_shuffle[6336];
    assign key_original[2652] = key_shuffle[1917];
    assign key_original[2651] = key_shuffle[7057];
    assign key_original[2650] = key_shuffle[3278];
    assign key_original[2649] = key_shuffle[6611];
    assign key_original[2648] = key_shuffle[7925];
    assign key_original[2647] = key_shuffle[2931];
    assign key_original[2646] = key_shuffle[6434];
    assign key_original[2645] = key_shuffle[8160];
    assign key_original[2644] = key_shuffle[4548];
    assign key_original[2643] = key_shuffle[2425];
    assign key_original[2642] = key_shuffle[1828];
    assign key_original[2641] = key_shuffle[4322];
    assign key_original[2640] = key_shuffle[1805];
    assign key_original[2639] = key_shuffle[5487];
    assign key_original[2638] = key_shuffle[2847];
    assign key_original[2637] = key_shuffle[5862];
    assign key_original[2636] = key_shuffle[599];
    assign key_original[2635] = key_shuffle[7918];
    assign key_original[2634] = key_shuffle[7012];
    assign key_original[2633] = key_shuffle[3113];
    assign key_original[2632] = key_shuffle[1505];
    assign key_original[2631] = key_shuffle[3790];
    assign key_original[2630] = key_shuffle[2741];
    assign key_original[2629] = key_shuffle[363];
    assign key_original[2628] = key_shuffle[1445];
    assign key_original[2627] = key_shuffle[4466];
    assign key_original[2626] = key_shuffle[1082];
    assign key_original[2625] = key_shuffle[1930];
    assign key_original[2624] = key_shuffle[1529];
    assign key_original[2623] = key_shuffle[23];
    assign key_original[2622] = key_shuffle[2336];
    assign key_original[2621] = key_shuffle[1391];
    assign key_original[2620] = key_shuffle[6602];
    assign key_original[2619] = key_shuffle[5950];
    assign key_original[2618] = key_shuffle[5195];
    assign key_original[2617] = key_shuffle[6796];
    assign key_original[2616] = key_shuffle[4469];
    assign key_original[2615] = key_shuffle[5865];
    assign key_original[2614] = key_shuffle[5679];
    assign key_original[2613] = key_shuffle[7687];
    assign key_original[2612] = key_shuffle[5642];
    assign key_original[2611] = key_shuffle[6351];
    assign key_original[2610] = key_shuffle[7648];
    assign key_original[2609] = key_shuffle[1972];
    assign key_original[2608] = key_shuffle[7340];
    assign key_original[2607] = key_shuffle[4510];
    assign key_original[2606] = key_shuffle[4974];
    assign key_original[2605] = key_shuffle[7304];
    assign key_original[2604] = key_shuffle[3352];
    assign key_original[2603] = key_shuffle[3196];
    assign key_original[2602] = key_shuffle[3657];
    assign key_original[2601] = key_shuffle[4479];
    assign key_original[2600] = key_shuffle[7531];
    assign key_original[2599] = key_shuffle[6950];
    assign key_original[2598] = key_shuffle[4046];
    assign key_original[2597] = key_shuffle[4387];
    assign key_original[2596] = key_shuffle[2570];
    assign key_original[2595] = key_shuffle[5341];
    assign key_original[2594] = key_shuffle[5841];
    assign key_original[2593] = key_shuffle[5337];
    assign key_original[2592] = key_shuffle[6936];
    assign key_original[2591] = key_shuffle[4637];
    assign key_original[2590] = key_shuffle[8063];
    assign key_original[2589] = key_shuffle[360];
    assign key_original[2588] = key_shuffle[7289];
    assign key_original[2587] = key_shuffle[3566];
    assign key_original[2586] = key_shuffle[4798];
    assign key_original[2585] = key_shuffle[5535];
    assign key_original[2584] = key_shuffle[2178];
    assign key_original[2583] = key_shuffle[5152];
    assign key_original[2582] = key_shuffle[6111];
    assign key_original[2581] = key_shuffle[3005];
    assign key_original[2580] = key_shuffle[1896];
    assign key_original[2579] = key_shuffle[4044];
    assign key_original[2578] = key_shuffle[918];
    assign key_original[2577] = key_shuffle[5283];
    assign key_original[2576] = key_shuffle[7235];
    assign key_original[2575] = key_shuffle[607];
    assign key_original[2574] = key_shuffle[7183];
    assign key_original[2573] = key_shuffle[2001];
    assign key_original[2572] = key_shuffle[4982];
    assign key_original[2571] = key_shuffle[6892];
    assign key_original[2570] = key_shuffle[287];
    assign key_original[2569] = key_shuffle[4894];
    assign key_original[2568] = key_shuffle[6767];
    assign key_original[2567] = key_shuffle[7324];
    assign key_original[2566] = key_shuffle[4445];
    assign key_original[2565] = key_shuffle[950];
    assign key_original[2564] = key_shuffle[4562];
    assign key_original[2563] = key_shuffle[1604];
    assign key_original[2562] = key_shuffle[6664];
    assign key_original[2561] = key_shuffle[7936];
    assign key_original[2560] = key_shuffle[3227];
    assign key_original[2559] = key_shuffle[7921];
    assign key_original[2558] = key_shuffle[831];
    assign key_original[2557] = key_shuffle[5053];
    assign key_original[2556] = key_shuffle[7205];
    assign key_original[2555] = key_shuffle[7483];
    assign key_original[2554] = key_shuffle[6218];
    assign key_original[2553] = key_shuffle[6831];
    assign key_original[2552] = key_shuffle[7471];
    assign key_original[2551] = key_shuffle[4128];
    assign key_original[2550] = key_shuffle[232];
    assign key_original[2549] = key_shuffle[3845];
    assign key_original[2548] = key_shuffle[4772];
    assign key_original[2547] = key_shuffle[6942];
    assign key_original[2546] = key_shuffle[5458];
    assign key_original[2545] = key_shuffle[723];
    assign key_original[2544] = key_shuffle[3249];
    assign key_original[2543] = key_shuffle[6961];
    assign key_original[2542] = key_shuffle[6413];
    assign key_original[2541] = key_shuffle[8007];
    assign key_original[2540] = key_shuffle[1934];
    assign key_original[2539] = key_shuffle[6762];
    assign key_original[2538] = key_shuffle[2051];
    assign key_original[2537] = key_shuffle[5020];
    assign key_original[2536] = key_shuffle[405];
    assign key_original[2535] = key_shuffle[6778];
    assign key_original[2534] = key_shuffle[504];
    assign key_original[2533] = key_shuffle[7584];
    assign key_original[2532] = key_shuffle[5102];
    assign key_original[2531] = key_shuffle[6427];
    assign key_original[2530] = key_shuffle[501];
    assign key_original[2529] = key_shuffle[7418];
    assign key_original[2528] = key_shuffle[4985];
    assign key_original[2527] = key_shuffle[2066];
    assign key_original[2526] = key_shuffle[7933];
    assign key_original[2525] = key_shuffle[1885];
    assign key_original[2524] = key_shuffle[5762];
    assign key_original[2523] = key_shuffle[6735];
    assign key_original[2522] = key_shuffle[5946];
    assign key_original[2521] = key_shuffle[7106];
    assign key_original[2520] = key_shuffle[4860];
    assign key_original[2519] = key_shuffle[8166];
    assign key_original[2518] = key_shuffle[7279];
    assign key_original[2517] = key_shuffle[1157];
    assign key_original[2516] = key_shuffle[1443];
    assign key_original[2515] = key_shuffle[8109];
    assign key_original[2514] = key_shuffle[7769];
    assign key_original[2513] = key_shuffle[7136];
    assign key_original[2512] = key_shuffle[7440];
    assign key_original[2511] = key_shuffle[839];
    assign key_original[2510] = key_shuffle[521];
    assign key_original[2509] = key_shuffle[7162];
    assign key_original[2508] = key_shuffle[1297];
    assign key_original[2507] = key_shuffle[2194];
    assign key_original[2506] = key_shuffle[4432];
    assign key_original[2505] = key_shuffle[5128];
    assign key_original[2504] = key_shuffle[6065];
    assign key_original[2503] = key_shuffle[5765];
    assign key_original[2502] = key_shuffle[6790];
    assign key_original[2501] = key_shuffle[3757];
    assign key_original[2500] = key_shuffle[4471];
    assign key_original[2499] = key_shuffle[4225];
    assign key_original[2498] = key_shuffle[1605];
    assign key_original[2497] = key_shuffle[4035];
    assign key_original[2496] = key_shuffle[6545];
    assign key_original[2495] = key_shuffle[7892];
    assign key_original[2494] = key_shuffle[2322];
    assign key_original[2493] = key_shuffle[7227];
    assign key_original[2492] = key_shuffle[7672];
    assign key_original[2491] = key_shuffle[6630];
    assign key_original[2490] = key_shuffle[6937];
    assign key_original[2489] = key_shuffle[2796];
    assign key_original[2488] = key_shuffle[525];
    assign key_original[2487] = key_shuffle[6491];
    assign key_original[2486] = key_shuffle[3980];
    assign key_original[2485] = key_shuffle[2529];
    assign key_original[2484] = key_shuffle[3848];
    assign key_original[2483] = key_shuffle[4849];
    assign key_original[2482] = key_shuffle[2146];
    assign key_original[2481] = key_shuffle[6988];
    assign key_original[2480] = key_shuffle[5094];
    assign key_original[2479] = key_shuffle[4865];
    assign key_original[2478] = key_shuffle[2215];
    assign key_original[2477] = key_shuffle[7560];
    assign key_original[2476] = key_shuffle[3737];
    assign key_original[2475] = key_shuffle[5205];
    assign key_original[2474] = key_shuffle[5079];
    assign key_original[2473] = key_shuffle[1810];
    assign key_original[2472] = key_shuffle[4862];
    assign key_original[2471] = key_shuffle[1501];
    assign key_original[2470] = key_shuffle[7408];
    assign key_original[2469] = key_shuffle[5611];
    assign key_original[2468] = key_shuffle[3242];
    assign key_original[2467] = key_shuffle[5445];
    assign key_original[2466] = key_shuffle[264];
    assign key_original[2465] = key_shuffle[2655];
    assign key_original[2464] = key_shuffle[6236];
    assign key_original[2463] = key_shuffle[2299];
    assign key_original[2462] = key_shuffle[1516];
    assign key_original[2461] = key_shuffle[61];
    assign key_original[2460] = key_shuffle[4613];
    assign key_original[2459] = key_shuffle[1255];
    assign key_original[2458] = key_shuffle[3319];
    assign key_original[2457] = key_shuffle[6490];
    assign key_original[2456] = key_shuffle[1781];
    assign key_original[2455] = key_shuffle[6326];
    assign key_original[2454] = key_shuffle[484];
    assign key_original[2453] = key_shuffle[6105];
    assign key_original[2452] = key_shuffle[7840];
    assign key_original[2451] = key_shuffle[1770];
    assign key_original[2450] = key_shuffle[5014];
    assign key_original[2449] = key_shuffle[7545];
    assign key_original[2448] = key_shuffle[6895];
    assign key_original[2447] = key_shuffle[6614];
    assign key_original[2446] = key_shuffle[5842];
    assign key_original[2445] = key_shuffle[897];
    assign key_original[2444] = key_shuffle[5722];
    assign key_original[2443] = key_shuffle[6751];
    assign key_original[2442] = key_shuffle[1122];
    assign key_original[2441] = key_shuffle[6764];
    assign key_original[2440] = key_shuffle[6188];
    assign key_original[2439] = key_shuffle[675];
    assign key_original[2438] = key_shuffle[4184];
    assign key_original[2437] = key_shuffle[4365];
    assign key_original[2436] = key_shuffle[3713];
    assign key_original[2435] = key_shuffle[2970];
    assign key_original[2434] = key_shuffle[637];
    assign key_original[2433] = key_shuffle[252];
    assign key_original[2432] = key_shuffle[1656];
    assign key_original[2431] = key_shuffle[4165];
    assign key_original[2430] = key_shuffle[3764];
    assign key_original[2429] = key_shuffle[7688];
    assign key_original[2428] = key_shuffle[6514];
    assign key_original[2427] = key_shuffle[489];
    assign key_original[2426] = key_shuffle[2067];
    assign key_original[2425] = key_shuffle[2573];
    assign key_original[2424] = key_shuffle[7573];
    assign key_original[2423] = key_shuffle[767];
    assign key_original[2422] = key_shuffle[5531];
    assign key_original[2421] = key_shuffle[1666];
    assign key_original[2420] = key_shuffle[3507];
    assign key_original[2419] = key_shuffle[5247];
    assign key_original[2418] = key_shuffle[999];
    assign key_original[2417] = key_shuffle[568];
    assign key_original[2416] = key_shuffle[1264];
    assign key_original[2415] = key_shuffle[33];
    assign key_original[2414] = key_shuffle[6143];
    assign key_original[2413] = key_shuffle[4820];
    assign key_original[2412] = key_shuffle[2330];
    assign key_original[2411] = key_shuffle[8070];
    assign key_original[2410] = key_shuffle[2449];
    assign key_original[2409] = key_shuffle[7041];
    assign key_original[2408] = key_shuffle[7058];
    assign key_original[2407] = key_shuffle[5621];
    assign key_original[2406] = key_shuffle[2131];
    assign key_original[2405] = key_shuffle[1655];
    assign key_original[2404] = key_shuffle[257];
    assign key_original[2403] = key_shuffle[1373];
    assign key_original[2402] = key_shuffle[4715];
    assign key_original[2401] = key_shuffle[6609];
    assign key_original[2400] = key_shuffle[8066];
    assign key_original[2399] = key_shuffle[2361];
    assign key_original[2398] = key_shuffle[4358];
    assign key_original[2397] = key_shuffle[7820];
    assign key_original[2396] = key_shuffle[6070];
    assign key_original[2395] = key_shuffle[3431];
    assign key_original[2394] = key_shuffle[4367];
    assign key_original[2393] = key_shuffle[6619];
    assign key_original[2392] = key_shuffle[5798];
    assign key_original[2391] = key_shuffle[7220];
    assign key_original[2390] = key_shuffle[1569];
    assign key_original[2389] = key_shuffle[361];
    assign key_original[2388] = key_shuffle[366];
    assign key_original[2387] = key_shuffle[2617];
    assign key_original[2386] = key_shuffle[7745];
    assign key_original[2385] = key_shuffle[7765];
    assign key_original[2384] = key_shuffle[3360];
    assign key_original[2383] = key_shuffle[6595];
    assign key_original[2382] = key_shuffle[1916];
    assign key_original[2381] = key_shuffle[2484];
    assign key_original[2380] = key_shuffle[5273];
    assign key_original[2379] = key_shuffle[2468];
    assign key_original[2378] = key_shuffle[267];
    assign key_original[2377] = key_shuffle[1554];
    assign key_original[2376] = key_shuffle[211];
    assign key_original[2375] = key_shuffle[7863];
    assign key_original[2374] = key_shuffle[8183];
    assign key_original[2373] = key_shuffle[887];
    assign key_original[2372] = key_shuffle[1313];
    assign key_original[2371] = key_shuffle[3988];
    assign key_original[2370] = key_shuffle[1820];
    assign key_original[2369] = key_shuffle[2384];
    assign key_original[2368] = key_shuffle[7318];
    assign key_original[2367] = key_shuffle[5709];
    assign key_original[2366] = key_shuffle[3948];
    assign key_original[2365] = key_shuffle[154];
    assign key_original[2364] = key_shuffle[5756];
    assign key_original[2363] = key_shuffle[4072];
    assign key_original[2362] = key_shuffle[1578];
    assign key_original[2361] = key_shuffle[2936];
    assign key_original[2360] = key_shuffle[1707];
    assign key_original[2359] = key_shuffle[4130];
    assign key_original[2358] = key_shuffle[4085];
    assign key_original[2357] = key_shuffle[3674];
    assign key_original[2356] = key_shuffle[5356];
    assign key_original[2355] = key_shuffle[6774];
    assign key_original[2354] = key_shuffle[101];
    assign key_original[2353] = key_shuffle[648];
    assign key_original[2352] = key_shuffle[384];
    assign key_original[2351] = key_shuffle[694];
    assign key_original[2350] = key_shuffle[369];
    assign key_original[2349] = key_shuffle[2709];
    assign key_original[2348] = key_shuffle[1937];
    assign key_original[2347] = key_shuffle[4107];
    assign key_original[2346] = key_shuffle[3415];
    assign key_original[2345] = key_shuffle[8000];
    assign key_original[2344] = key_shuffle[994];
    assign key_original[2343] = key_shuffle[2625];
    assign key_original[2342] = key_shuffle[5799];
    assign key_original[2341] = key_shuffle[4106];
    assign key_original[2340] = key_shuffle[4401];
    assign key_original[2339] = key_shuffle[5335];
    assign key_original[2338] = key_shuffle[4301];
    assign key_original[2337] = key_shuffle[5293];
    assign key_original[2336] = key_shuffle[3896];
    assign key_original[2335] = key_shuffle[263];
    assign key_original[2334] = key_shuffle[2800];
    assign key_original[2333] = key_shuffle[2972];
    assign key_original[2332] = key_shuffle[3585];
    assign key_original[2331] = key_shuffle[1513];
    assign key_original[2330] = key_shuffle[6907];
    assign key_original[2329] = key_shuffle[7438];
    assign key_original[2328] = key_shuffle[6181];
    assign key_original[2327] = key_shuffle[498];
    assign key_original[2326] = key_shuffle[153];
    assign key_original[2325] = key_shuffle[6674];
    assign key_original[2324] = key_shuffle[2722];
    assign key_original[2323] = key_shuffle[7007];
    assign key_original[2322] = key_shuffle[906];
    assign key_original[2321] = key_shuffle[4381];
    assign key_original[2320] = key_shuffle[5193];
    assign key_original[2319] = key_shuffle[4895];
    assign key_original[2318] = key_shuffle[1508];
    assign key_original[2317] = key_shuffle[6061];
    assign key_original[2316] = key_shuffle[3111];
    assign key_original[2315] = key_shuffle[548];
    assign key_original[2314] = key_shuffle[5395];
    assign key_original[2313] = key_shuffle[7109];
    assign key_original[2312] = key_shuffle[6945];
    assign key_original[2311] = key_shuffle[1193];
    assign key_original[2310] = key_shuffle[5580];
    assign key_original[2309] = key_shuffle[6931];
    assign key_original[2308] = key_shuffle[4482];
    assign key_original[2307] = key_shuffle[1198];
    assign key_original[2306] = key_shuffle[5781];
    assign key_original[2305] = key_shuffle[6893];
    assign key_original[2304] = key_shuffle[5991];
    assign key_original[2303] = key_shuffle[1403];
    assign key_original[2302] = key_shuffle[2495];
    assign key_original[2301] = key_shuffle[2164];
    assign key_original[2300] = key_shuffle[3808];
    assign key_original[2299] = key_shuffle[7827];
    assign key_original[2298] = key_shuffle[4929];
    assign key_original[2297] = key_shuffle[3554];
    assign key_original[2296] = key_shuffle[5180];
    assign key_original[2295] = key_shuffle[5966];
    assign key_original[2294] = key_shuffle[6891];
    assign key_original[2293] = key_shuffle[4903];
    assign key_original[2292] = key_shuffle[4949];
    assign key_original[2291] = key_shuffle[1208];
    assign key_original[2290] = key_shuffle[5868];
    assign key_original[2289] = key_shuffle[6148];
    assign key_original[2288] = key_shuffle[3018];
    assign key_original[2287] = key_shuffle[870];
    assign key_original[2286] = key_shuffle[1690];
    assign key_original[2285] = key_shuffle[7977];
    assign key_original[2284] = key_shuffle[5384];
    assign key_original[2283] = key_shuffle[2943];
    assign key_original[2282] = key_shuffle[7363];
    assign key_original[2281] = key_shuffle[4450];
    assign key_original[2280] = key_shuffle[2317];
    assign key_original[2279] = key_shuffle[6443];
    assign key_original[2278] = key_shuffle[6482];
    assign key_original[2277] = key_shuffle[1155];
    assign key_original[2276] = key_shuffle[128];
    assign key_original[2275] = key_shuffle[5931];
    assign key_original[2274] = key_shuffle[3716];
    assign key_original[2273] = key_shuffle[7662];
    assign key_original[2272] = key_shuffle[7285];
    assign key_original[2271] = key_shuffle[895];
    assign key_original[2270] = key_shuffle[7457];
    assign key_original[2269] = key_shuffle[3999];
    assign key_original[2268] = key_shuffle[2864];
    assign key_original[2267] = key_shuffle[6519];
    assign key_original[2266] = key_shuffle[3583];
    assign key_original[2265] = key_shuffle[454];
    assign key_original[2264] = key_shuffle[54];
    assign key_original[2263] = key_shuffle[6526];
    assign key_original[2262] = key_shuffle[2777];
    assign key_original[2261] = key_shuffle[5499];
    assign key_original[2260] = key_shuffle[1027];
    assign key_original[2259] = key_shuffle[3006];
    assign key_original[2258] = key_shuffle[505];
    assign key_original[2257] = key_shuffle[6858];
    assign key_original[2256] = key_shuffle[3899];
    assign key_original[2255] = key_shuffle[3637];
    assign key_original[2254] = key_shuffle[5342];
    assign key_original[2253] = key_shuffle[1435];
    assign key_original[2252] = key_shuffle[4018];
    assign key_original[2251] = key_shuffle[5929];
    assign key_original[2250] = key_shuffle[7053];
    assign key_original[2249] = key_shuffle[793];
    assign key_original[2248] = key_shuffle[6620];
    assign key_original[2247] = key_shuffle[3871];
    assign key_original[2246] = key_shuffle[4066];
    assign key_original[2245] = key_shuffle[3650];
    assign key_original[2244] = key_shuffle[49];
    assign key_original[2243] = key_shuffle[1822];
    assign key_original[2242] = key_shuffle[2103];
    assign key_original[2241] = key_shuffle[2086];
    assign key_original[2240] = key_shuffle[6076];
    assign key_original[2239] = key_shuffle[589];
    assign key_original[2238] = key_shuffle[8145];
    assign key_original[2237] = key_shuffle[6064];
    assign key_original[2236] = key_shuffle[8060];
    assign key_original[2235] = key_shuffle[4529];
    assign key_original[2234] = key_shuffle[5596];
    assign key_original[2233] = key_shuffle[5114];
    assign key_original[2232] = key_shuffle[1977];
    assign key_original[2231] = key_shuffle[3917];
    assign key_original[2230] = key_shuffle[4742];
    assign key_original[2229] = key_shuffle[2415];
    assign key_original[2228] = key_shuffle[6437];
    assign key_original[2227] = key_shuffle[8125];
    assign key_original[2226] = key_shuffle[6784];
    assign key_original[2225] = key_shuffle[4959];
    assign key_original[2224] = key_shuffle[1274];
    assign key_original[2223] = key_shuffle[3357];
    assign key_original[2222] = key_shuffle[3557];
    assign key_original[2221] = key_shuffle[5430];
    assign key_original[2220] = key_shuffle[1665];
    assign key_original[2219] = key_shuffle[3959];
    assign key_original[2218] = key_shuffle[4242];
    assign key_original[2217] = key_shuffle[1309];
    assign key_original[2216] = key_shuffle[3789];
    assign key_original[2215] = key_shuffle[2990];
    assign key_original[2214] = key_shuffle[846];
    assign key_original[2213] = key_shuffle[3230];
    assign key_original[2212] = key_shuffle[142];
    assign key_original[2211] = key_shuffle[6023];
    assign key_original[2210] = key_shuffle[4235];
    assign key_original[2209] = key_shuffle[3593];
    assign key_original[2208] = key_shuffle[6706];
    assign key_original[2207] = key_shuffle[784];
    assign key_original[2206] = key_shuffle[3039];
    assign key_original[2205] = key_shuffle[5112];
    assign key_original[2204] = key_shuffle[4736];
    assign key_original[2203] = key_shuffle[4571];
    assign key_original[2202] = key_shuffle[986];
    assign key_original[2201] = key_shuffle[1565];
    assign key_original[2200] = key_shuffle[7277];
    assign key_original[2199] = key_shuffle[50];
    assign key_original[2198] = key_shuffle[6327];
    assign key_original[2197] = key_shuffle[3575];
    assign key_original[2196] = key_shuffle[7740];
    assign key_original[2195] = key_shuffle[452];
    assign key_original[2194] = key_shuffle[6320];
    assign key_original[2193] = key_shuffle[1076];
    assign key_original[2192] = key_shuffle[799];
    assign key_original[2191] = key_shuffle[4528];
    assign key_original[2190] = key_shuffle[2133];
    assign key_original[2189] = key_shuffle[3887];
    assign key_original[2188] = key_shuffle[7492];
    assign key_original[2187] = key_shuffle[5554];
    assign key_original[2186] = key_shuffle[5457];
    assign key_original[2185] = key_shuffle[4976];
    assign key_original[2184] = key_shuffle[1796];
    assign key_original[2183] = key_shuffle[6008];
    assign key_original[2182] = key_shuffle[2889];
    assign key_original[2181] = key_shuffle[6400];
    assign key_original[2180] = key_shuffle[1658];
    assign key_original[2179] = key_shuffle[5790];
    assign key_original[2178] = key_shuffle[2225];
    assign key_original[2177] = key_shuffle[1244];
    assign key_original[2176] = key_shuffle[6321];
    assign key_original[2175] = key_shuffle[2243];
    assign key_original[2174] = key_shuffle[3533];
    assign key_original[2173] = key_shuffle[6569];
    assign key_original[2172] = key_shuffle[3571];
    assign key_original[2171] = key_shuffle[5586];
    assign key_original[2170] = key_shuffle[6965];
    assign key_original[2169] = key_shuffle[4832];
    assign key_original[2168] = key_shuffle[2020];
    assign key_original[2167] = key_shuffle[2070];
    assign key_original[2166] = key_shuffle[1778];
    assign key_original[2165] = key_shuffle[14];
    assign key_original[2164] = key_shuffle[7610];
    assign key_original[2163] = key_shuffle[3069];
    assign key_original[2162] = key_shuffle[4618];
    assign key_original[2161] = key_shuffle[5416];
    assign key_original[2160] = key_shuffle[1194];
    assign key_original[2159] = key_shuffle[4504];
    assign key_original[2158] = key_shuffle[5423];
    assign key_original[2157] = key_shuffle[562];
    assign key_original[2156] = key_shuffle[4789];
    assign key_original[2155] = key_shuffle[341];
    assign key_original[2154] = key_shuffle[5407];
    assign key_original[2153] = key_shuffle[6703];
    assign key_original[2152] = key_shuffle[4374];
    assign key_original[2151] = key_shuffle[4098];
    assign key_original[2150] = key_shuffle[6050];
    assign key_original[2149] = key_shuffle[4443];
    assign key_original[2148] = key_shuffle[5987];
    assign key_original[2147] = key_shuffle[843];
    assign key_original[2146] = key_shuffle[5204];
    assign key_original[2145] = key_shuffle[1682];
    assign key_original[2144] = key_shuffle[6441];
    assign key_original[2143] = key_shuffle[7917];
    assign key_original[2142] = key_shuffle[7138];
    assign key_original[2141] = key_shuffle[995];
    assign key_original[2140] = key_shuffle[5133];
    assign key_original[2139] = key_shuffle[7249];
    assign key_original[2138] = key_shuffle[7474];
    assign key_original[2137] = key_shuffle[4245];
    assign key_original[2136] = key_shuffle[2395];
    assign key_original[2135] = key_shuffle[2761];
    assign key_original[2134] = key_shuffle[5137];
    assign key_original[2133] = key_shuffle[6080];
    assign key_original[2132] = key_shuffle[5403];
    assign key_original[2131] = key_shuffle[6041];
    assign key_original[2130] = key_shuffle[4102];
    assign key_original[2129] = key_shuffle[1436];
    assign key_original[2128] = key_shuffle[2237];
    assign key_original[2127] = key_shuffle[8126];
    assign key_original[2126] = key_shuffle[1050];
    assign key_original[2125] = key_shuffle[4899];
    assign key_original[2124] = key_shuffle[5849];
    assign key_original[2123] = key_shuffle[91];
    assign key_original[2122] = key_shuffle[1067];
    assign key_original[2121] = key_shuffle[960];
    assign key_original[2120] = key_shuffle[537];
    assign key_original[2119] = key_shuffle[4752];
    assign key_original[2118] = key_shuffle[1095];
    assign key_original[2117] = key_shuffle[6135];
    assign key_original[2116] = key_shuffle[446];
    assign key_original[2115] = key_shuffle[6486];
    assign key_original[2114] = key_shuffle[759];
    assign key_original[2113] = key_shuffle[6110];
    assign key_original[2112] = key_shuffle[7524];
    assign key_original[2111] = key_shuffle[526];
    assign key_original[2110] = key_shuffle[6849];
    assign key_original[2109] = key_shuffle[4735];
    assign key_original[2108] = key_shuffle[320];
    assign key_original[2107] = key_shuffle[2868];
    assign key_original[2106] = key_shuffle[3804];
    assign key_original[2105] = key_shuffle[6828];
    assign key_original[2104] = key_shuffle[6275];
    assign key_original[2103] = key_shuffle[2142];
    assign key_original[2102] = key_shuffle[7431];
    assign key_original[2101] = key_shuffle[766];
    assign key_original[2100] = key_shuffle[7286];
    assign key_original[2099] = key_shuffle[355];
    assign key_original[2098] = key_shuffle[1123];
    assign key_original[2097] = key_shuffle[5900];
    assign key_original[2096] = key_shuffle[1976];
    assign key_original[2095] = key_shuffle[3924];
    assign key_original[2094] = key_shuffle[5810];
    assign key_original[2093] = key_shuffle[2974];
    assign key_original[2092] = key_shuffle[5368];
    assign key_original[2091] = key_shuffle[2921];
    assign key_original[2090] = key_shuffle[7021];
    assign key_original[2089] = key_shuffle[2467];
    assign key_original[2088] = key_shuffle[7758];
    assign key_original[2087] = key_shuffle[4139];
    assign key_original[2086] = key_shuffle[4131];
    assign key_original[2085] = key_shuffle[6991];
    assign key_original[2084] = key_shuffle[6027];
    assign key_original[2083] = key_shuffle[6547];
    assign key_original[2082] = key_shuffle[4629];
    assign key_original[2081] = key_shuffle[5983];
    assign key_original[2080] = key_shuffle[476];
    assign key_original[2079] = key_shuffle[6485];
    assign key_original[2078] = key_shuffle[2618];
    assign key_original[2077] = key_shuffle[284];
    assign key_original[2076] = key_shuffle[6253];
    assign key_original[2075] = key_shuffle[810];
    assign key_original[2074] = key_shuffle[883];
    assign key_original[2073] = key_shuffle[7081];
    assign key_original[2072] = key_shuffle[2473];
    assign key_original[2071] = key_shuffle[3981];
    assign key_original[2070] = key_shuffle[3517];
    assign key_original[2069] = key_shuffle[6742];
    assign key_original[2068] = key_shuffle[1661];
    assign key_original[2067] = key_shuffle[2239];
    assign key_original[2066] = key_shuffle[5662];
    assign key_original[2065] = key_shuffle[7132];
    assign key_original[2064] = key_shuffle[4604];
    assign key_original[2063] = key_shuffle[3264];
    assign key_original[2062] = key_shuffle[4160];
    assign key_original[2061] = key_shuffle[8019];
    assign key_original[2060] = key_shuffle[5825];
    assign key_original[2059] = key_shuffle[6391];
    assign key_original[2058] = key_shuffle[3321];
    assign key_original[2057] = key_shuffle[4680];
    assign key_original[2056] = key_shuffle[3581];
    assign key_original[2055] = key_shuffle[673];
    assign key_original[2054] = key_shuffle[7365];
    assign key_original[2053] = key_shuffle[2826];
    assign key_original[2052] = key_shuffle[5131];
    assign key_original[2051] = key_shuffle[6698];
    assign key_original[2050] = key_shuffle[6675];
    assign key_original[2049] = key_shuffle[3691];
    assign key_original[2048] = key_shuffle[5129];
    assign key_original[2047] = key_shuffle[5904];
    assign key_original[2046] = key_shuffle[6260];
    assign key_original[2045] = key_shuffle[7215];
    assign key_original[2044] = key_shuffle[7060];
    assign key_original[2043] = key_shuffle[559];
    assign key_original[2042] = key_shuffle[2566];
    assign key_original[2041] = key_shuffle[7982];
    assign key_original[2040] = key_shuffle[2226];
    assign key_original[2039] = key_shuffle[4483];
    assign key_original[2038] = key_shuffle[7209];
    assign key_original[2037] = key_shuffle[1001];
    assign key_original[2036] = key_shuffle[7943];
    assign key_original[2035] = key_shuffle[262];
    assign key_original[2034] = key_shuffle[6466];
    assign key_original[2033] = key_shuffle[4439];
    assign key_original[2032] = key_shuffle[4697];
    assign key_original[2031] = key_shuffle[3596];
    assign key_original[2030] = key_shuffle[1973];
    assign key_original[2029] = key_shuffle[777];
    assign key_original[2028] = key_shuffle[84];
    assign key_original[2027] = key_shuffle[3488];
    assign key_original[2026] = key_shuffle[1939];
    assign key_original[2025] = key_shuffle[1110];
    assign key_original[2024] = key_shuffle[4038];
    assign key_original[2023] = key_shuffle[2496];
    assign key_original[2022] = key_shuffle[6460];
    assign key_original[2021] = key_shuffle[6368];
    assign key_original[2020] = key_shuffle[4666];
    assign key_original[2019] = key_shuffle[4705];
    assign key_original[2018] = key_shuffle[3992];
    assign key_original[2017] = key_shuffle[4864];
    assign key_original[2016] = key_shuffle[908];
    assign key_original[2015] = key_shuffle[6914];
    assign key_original[2014] = key_shuffle[4769];
    assign key_original[2013] = key_shuffle[6383];
    assign key_original[2012] = key_shuffle[5906];
    assign key_original[2011] = key_shuffle[5396];
    assign key_original[2010] = key_shuffle[7851];
    assign key_original[2009] = key_shuffle[6865];
    assign key_original[2008] = key_shuffle[5387];
    assign key_original[2007] = key_shuffle[642];
    assign key_original[2006] = key_shuffle[4061];
    assign key_original[2005] = key_shuffle[1412];
    assign key_original[2004] = key_shuffle[4563];
    assign key_original[2003] = key_shuffle[7913];
    assign key_original[2002] = key_shuffle[5704];
    assign key_original[2001] = key_shuffle[497];
    assign key_original[2000] = key_shuffle[1481];
    assign key_original[1999] = key_shuffle[2478];
    assign key_original[1998] = key_shuffle[7201];
    assign key_original[1997] = key_shuffle[5763];
    assign key_original[1996] = key_shuffle[2159];
    assign key_original[1995] = key_shuffle[6082];
    assign key_original[1994] = key_shuffle[7236];
    assign key_original[1993] = key_shuffle[1620];
    assign key_original[1992] = key_shuffle[5272];
    assign key_original[1991] = key_shuffle[7633];
    assign key_original[1990] = key_shuffle[2592];
    assign key_original[1989] = key_shuffle[2165];
    assign key_original[1988] = key_shuffle[4083];
    assign key_original[1987] = key_shuffle[6806];
    assign key_original[1986] = key_shuffle[3736];
    assign key_original[1985] = key_shuffle[6660];
    assign key_original[1984] = key_shuffle[3686];
    assign key_original[1983] = key_shuffle[6911];
    assign key_original[1982] = key_shuffle[2362];
    assign key_original[1981] = key_shuffle[886];
    assign key_original[1980] = key_shuffle[3330];
    assign key_original[1979] = key_shuffle[3562];
    assign key_original[1978] = key_shuffle[2244];
    assign key_original[1977] = key_shuffle[4191];
    assign key_original[1976] = key_shuffle[7185];
    assign key_original[1975] = key_shuffle[6736];
    assign key_original[1974] = key_shuffle[253];
    assign key_original[1973] = key_shuffle[7339];
    assign key_original[1972] = key_shuffle[7658];
    assign key_original[1971] = key_shuffle[8138];
    assign key_original[1970] = key_shuffle[4127];
    assign key_original[1969] = key_shuffle[5493];
    assign key_original[1968] = key_shuffle[2942];
    assign key_original[1967] = key_shuffle[2044];
    assign key_original[1966] = key_shuffle[5140];
    assign key_original[1965] = key_shuffle[2456];
    assign key_original[1964] = key_shuffle[5537];
    assign key_original[1963] = key_shuffle[68];
    assign key_original[1962] = key_shuffle[3485];
    assign key_original[1961] = key_shuffle[16];
    assign key_original[1960] = key_shuffle[4902];
    assign key_original[1959] = key_shuffle[978];
    assign key_original[1958] = key_shuffle[7655];
    assign key_original[1957] = key_shuffle[4186];
    assign key_original[1956] = key_shuffle[3704];
    assign key_original[1955] = key_shuffle[3292];
    assign key_original[1954] = key_shuffle[4656];
    assign key_original[1953] = key_shuffle[5192];
    assign key_original[1952] = key_shuffle[7487];
    assign key_original[1951] = key_shuffle[2364];
    assign key_original[1950] = key_shuffle[450];
    assign key_original[1949] = key_shuffle[2352];
    assign key_original[1948] = key_shuffle[5542];
    assign key_original[1947] = key_shuffle[5039];
    assign key_original[1946] = key_shuffle[1567];
    assign key_original[1945] = key_shuffle[7778];
    assign key_original[1944] = key_shuffle[3383];
    assign key_original[1943] = key_shuffle[7502];
    assign key_original[1942] = key_shuffle[5793];
    assign key_original[1941] = key_shuffle[4589];
    assign key_original[1940] = key_shuffle[4503];
    assign key_original[1939] = key_shuffle[2489];
    assign key_original[1938] = key_shuffle[685];
    assign key_original[1937] = key_shuffle[7099];
    assign key_original[1936] = key_shuffle[6913];
    assign key_original[1935] = key_shuffle[2650];
    assign key_original[1934] = key_shuffle[6101];
    assign key_original[1933] = key_shuffle[1572];
    assign key_original[1932] = key_shuffle[6415];
    assign key_original[1931] = key_shuffle[2409];
    assign key_original[1930] = key_shuffle[8164];
    assign key_original[1929] = key_shuffle[800];
    assign key_original[1928] = key_shuffle[6060];
    assign key_original[1927] = key_shuffle[281];
    assign key_original[1926] = key_shuffle[7629];
    assign key_original[1925] = key_shuffle[6948];
    assign key_original[1924] = key_shuffle[1135];
    assign key_original[1923] = key_shuffle[6337];
    assign key_original[1922] = key_shuffle[388];
    assign key_original[1921] = key_shuffle[32];
    assign key_original[1920] = key_shuffle[4868];
    assign key_original[1919] = key_shuffle[2094];
    assign key_original[1918] = key_shuffle[2038];
    assign key_original[1917] = key_shuffle[2869];
    assign key_original[1916] = key_shuffle[2134];
    assign key_original[1915] = key_shuffle[5447];
    assign key_original[1914] = key_shuffle[1696];
    assign key_original[1913] = key_shuffle[6395];
    assign key_original[1912] = key_shuffle[2753];
    assign key_original[1911] = key_shuffle[6740];
    assign key_original[1910] = key_shuffle[5489];
    assign key_original[1909] = key_shuffle[323];
    assign key_original[1908] = key_shuffle[5629];
    assign key_original[1907] = key_shuffle[4667];
    assign key_original[1906] = key_shuffle[6237];
    assign key_original[1905] = key_shuffle[6304];
    assign key_original[1904] = key_shuffle[1490];
    assign key_original[1903] = key_shuffle[7454];
    assign key_original[1902] = key_shuffle[3123];
    assign key_original[1901] = key_shuffle[4747];
    assign key_original[1900] = key_shuffle[2283];
    assign key_original[1899] = key_shuffle[5358];
    assign key_original[1898] = key_shuffle[7479];
    assign key_original[1897] = key_shuffle[6435];
    assign key_original[1896] = key_shuffle[4476];
    assign key_original[1895] = key_shuffle[737];
    assign key_original[1894] = key_shuffle[7384];
    assign key_original[1893] = key_shuffle[6507];
    assign key_original[1892] = key_shuffle[3873];
    assign key_original[1891] = key_shuffle[2746];
    assign key_original[1890] = key_shuffle[5869];
    assign key_original[1889] = key_shuffle[255];
    assign key_original[1888] = key_shuffle[1449];
    assign key_original[1887] = key_shuffle[2236];
    assign key_original[1886] = key_shuffle[2788];
    assign key_original[1885] = key_shuffle[3772];
    assign key_original[1884] = key_shuffle[5439];
    assign key_original[1883] = key_shuffle[1029];
    assign key_original[1882] = key_shuffle[6149];
    assign key_original[1881] = key_shuffle[300];
    assign key_original[1880] = key_shuffle[1310];
    assign key_original[1879] = key_shuffle[3903];
    assign key_original[1878] = key_shuffle[5072];
    assign key_original[1877] = key_shuffle[8034];
    assign key_original[1876] = key_shuffle[2170];
    assign key_original[1875] = key_shuffle[3475];
    assign key_original[1874] = key_shuffle[190];
    assign key_original[1873] = key_shuffle[606];
    assign key_original[1872] = key_shuffle[1447];
    assign key_original[1871] = key_shuffle[7239];
    assign key_original[1870] = key_shuffle[3240];
    assign key_original[1869] = key_shuffle[3774];
    assign key_original[1868] = key_shuffle[1108];
    assign key_original[1867] = key_shuffle[7577];
    assign key_original[1866] = key_shuffle[5209];
    assign key_original[1865] = key_shuffle[1068];
    assign key_original[1864] = key_shuffle[1823];
    assign key_original[1863] = key_shuffle[6283];
    assign key_original[1862] = key_shuffle[1575];
    assign key_original[1861] = key_shuffle[2917];
    assign key_original[1860] = key_shuffle[6870];
    assign key_original[1859] = key_shuffle[3487];
    assign key_original[1858] = key_shuffle[470];
    assign key_original[1857] = key_shuffle[7452];
    assign key_original[1856] = key_shuffle[275];
    assign key_original[1855] = key_shuffle[5646];
    assign key_original[1854] = key_shuffle[2181];
    assign key_original[1853] = key_shuffle[3798];
    assign key_original[1852] = key_shuffle[7467];
    assign key_original[1851] = key_shuffle[7412];
    assign key_original[1850] = key_shuffle[523];
    assign key_original[1849] = key_shuffle[2116];
    assign key_original[1848] = key_shuffle[3744];
    assign key_original[1847] = key_shuffle[4060];
    assign key_original[1846] = key_shuffle[6012];
    assign key_original[1845] = key_shuffle[7462];
    assign key_original[1844] = key_shuffle[5187];
    assign key_original[1843] = key_shuffle[1250];
    assign key_original[1842] = key_shuffle[770];
    assign key_original[1841] = key_shuffle[7341];
    assign key_original[1840] = key_shuffle[712];
    assign key_original[1839] = key_shuffle[4080];
    assign key_original[1838] = key_shuffle[1878];
    assign key_original[1837] = key_shuffle[7682];
    assign key_original[1836] = key_shuffle[2666];
    assign key_original[1835] = key_shuffle[6717];
    assign key_original[1834] = key_shuffle[2490];
    assign key_original[1833] = key_shuffle[4310];
    assign key_original[1832] = key_shuffle[3115];
    assign key_original[1831] = key_shuffle[3541];
    assign key_original[1830] = key_shuffle[2645];
    assign key_original[1829] = key_shuffle[2782];
    assign key_original[1828] = key_shuffle[582];
    assign key_original[1827] = key_shuffle[2046];
    assign key_original[1826] = key_shuffle[2144];
    assign key_original[1825] = key_shuffle[7311];
    assign key_original[1824] = key_shuffle[7754];
    assign key_original[1823] = key_shuffle[3291];
    assign key_original[1822] = key_shuffle[2772];
    assign key_original[1821] = key_shuffle[3432];
    assign key_original[1820] = key_shuffle[3679];
    assign key_original[1819] = key_shuffle[7383];
    assign key_original[1818] = key_shuffle[5155];
    assign key_original[1817] = key_shuffle[3695];
    assign key_original[1816] = key_shuffle[1777];
    assign key_original[1815] = key_shuffle[45];
    assign key_original[1814] = key_shuffle[3076];
    assign key_original[1813] = key_shuffle[969];
    assign key_original[1812] = key_shuffle[4135];
    assign key_original[1811] = key_shuffle[2379];
    assign key_original[1810] = key_shuffle[7693];
    assign key_original[1809] = key_shuffle[2844];
    assign key_original[1808] = key_shuffle[6940];
    assign key_original[1807] = key_shuffle[4920];
    assign key_original[1806] = key_shuffle[4525];
    assign key_original[1805] = key_shuffle[2270];
    assign key_original[1804] = key_shuffle[3694];
    assign key_original[1803] = key_shuffle[3690];
    assign key_original[1802] = key_shuffle[6031];
    assign key_original[1801] = key_shuffle[1214];
    assign key_original[1800] = key_shuffle[3205];
    assign key_original[1799] = key_shuffle[5113];
    assign key_original[1798] = key_shuffle[1348];
    assign key_original[1797] = key_shuffle[6886];
    assign key_original[1796] = key_shuffle[7419];
    assign key_original[1795] = key_shuffle[346];
    assign key_original[1794] = key_shuffle[6432];
    assign key_original[1793] = key_shuffle[5592];
    assign key_original[1792] = key_shuffle[4701];
    assign key_original[1791] = key_shuffle[2367];
    assign key_original[1790] = key_shuffle[7353];
    assign key_original[1789] = key_shuffle[7145];
    assign key_original[1788] = key_shuffle[1991];
    assign key_original[1787] = key_shuffle[5253];
    assign key_original[1786] = key_shuffle[4490];
    assign key_original[1785] = key_shuffle[1835];
    assign key_original[1784] = key_shuffle[5670];
    assign key_original[1783] = key_shuffle[6833];
    assign key_original[1782] = key_shuffle[4761];
    assign key_original[1781] = key_shuffle[2069];
    assign key_original[1780] = key_shuffle[3856];
    assign key_original[1779] = key_shuffle[4560];
    assign key_original[1778] = key_shuffle[216];
    assign key_original[1777] = key_shuffle[4379];
    assign key_original[1776] = key_shuffle[951];
    assign key_original[1775] = key_shuffle[3811];
    assign key_original[1774] = key_shuffle[1851];
    assign key_original[1773] = key_shuffle[1187];
    assign key_original[1772] = key_shuffle[7156];
    assign key_original[1771] = key_shuffle[2525];
    assign key_original[1770] = key_shuffle[433];
    assign key_original[1769] = key_shuffle[752];
    assign key_original[1768] = key_shuffle[7718];
    assign key_original[1767] = key_shuffle[103];
    assign key_original[1766] = key_shuffle[5139];
    assign key_original[1765] = key_shuffle[3519];
    assign key_original[1764] = key_shuffle[6976];
    assign key_original[1763] = key_shuffle[591];
    assign key_original[1762] = key_shuffle[6234];
    assign key_original[1761] = key_shuffle[6153];
    assign key_original[1760] = key_shuffle[5583];
    assign key_original[1759] = key_shuffle[6401];
    assign key_original[1758] = key_shuffle[2080];
    assign key_original[1757] = key_shuffle[4657];
    assign key_original[1756] = key_shuffle[605];
    assign key_original[1755] = key_shuffle[3800];
    assign key_original[1754] = key_shuffle[280];
    assign key_original[1753] = key_shuffle[4811];
    assign key_original[1752] = key_shuffle[6172];
    assign key_original[1751] = key_shuffle[6672];
    assign key_original[1750] = key_shuffle[2436];
    assign key_original[1749] = key_shuffle[5899];
    assign key_original[1748] = key_shuffle[7259];
    assign key_original[1747] = key_shuffle[1367];
    assign key_original[1746] = key_shuffle[6292];
    assign key_original[1745] = key_shuffle[1532];
    assign key_original[1744] = key_shuffle[4673];
    assign key_original[1743] = key_shuffle[2641];
    assign key_original[1742] = key_shuffle[1111];
    assign key_original[1741] = key_shuffle[6461];
    assign key_original[1740] = key_shuffle[2946];
    assign key_original[1739] = key_shuffle[842];
    assign key_original[1738] = key_shuffle[1455];
    assign key_original[1737] = key_shuffle[3652];
    assign key_original[1736] = key_shuffle[6267];
    assign key_original[1735] = key_shuffle[6433];
    assign key_original[1734] = key_shuffle[8061];
    assign key_original[1733] = key_shuffle[6568];
    assign key_original[1732] = key_shuffle[3163];
    assign key_original[1731] = key_shuffle[2639];
    assign key_original[1730] = key_shuffle[7118];
    assign key_original[1729] = key_shuffle[7026];
    assign key_original[1728] = key_shuffle[5672];
    assign key_original[1727] = key_shuffle[5286];
    assign key_original[1726] = key_shuffle[6097];
    assign key_original[1725] = key_shuffle[3553];
    assign key_original[1724] = key_shuffle[1697];
    assign key_original[1723] = key_shuffle[5323];
    assign key_original[1722] = key_shuffle[7589];
    assign key_original[1721] = key_shuffle[6637];
    assign key_original[1720] = key_shuffle[3200];
    assign key_original[1719] = key_shuffle[5059];
    assign key_original[1718] = key_shuffle[434];
    assign key_original[1717] = key_shuffle[3210];
    assign key_original[1716] = key_shuffle[3247];
    assign key_original[1715] = key_shuffle[5817];
    assign key_original[1714] = key_shuffle[8175];
    assign key_original[1713] = key_shuffle[1432];
    assign key_original[1712] = key_shuffle[2335];
    assign key_original[1711] = key_shuffle[7443];
    assign key_original[1710] = key_shuffle[2188];
    assign key_original[1709] = key_shuffle[5266];
    assign key_original[1708] = key_shuffle[3854];
    assign key_original[1707] = key_shuffle[3607];
    assign key_original[1706] = key_shuffle[3105];
    assign key_original[1705] = key_shuffle[4869];
    assign key_original[1704] = key_shuffle[6245];
    assign key_original[1703] = key_shuffle[1338];
    assign key_original[1702] = key_shuffle[3989];
    assign key_original[1701] = key_shuffle[7389];
    assign key_original[1700] = key_shuffle[7139];
    assign key_original[1699] = key_shuffle[1625];
    assign key_original[1698] = key_shuffle[3898];
    assign key_original[1697] = key_shuffle[5409];
    assign key_original[1696] = key_shuffle[7252];
    assign key_original[1695] = key_shuffle[4210];
    assign key_original[1694] = key_shuffle[4006];
    assign key_original[1693] = key_shuffle[909];
    assign key_original[1692] = key_shuffle[1594];
    assign key_original[1691] = key_shuffle[107];
    assign key_original[1690] = key_shuffle[2924];
    assign key_original[1689] = key_shuffle[4208];
    assign key_original[1688] = key_shuffle[2249];
    assign key_original[1687] = key_shuffle[3715];
    assign key_original[1686] = key_shuffle[528];
    assign key_original[1685] = key_shuffle[5243];
    assign key_original[1684] = key_shuffle[4318];
    assign key_original[1683] = key_shuffle[2346];
    assign key_original[1682] = key_shuffle[3429];
    assign key_original[1681] = key_shuffle[6623];
    assign key_original[1680] = key_shuffle[5319];
    assign key_original[1679] = key_shuffle[5644];
    assign key_original[1678] = key_shuffle[6373];
    assign key_original[1677] = key_shuffle[7051];
    assign key_original[1676] = key_shuffle[7518];
    assign key_original[1675] = key_shuffle[1000];
    assign key_original[1674] = key_shuffle[2672];
    assign key_original[1673] = key_shuffle[3970];
    assign key_original[1672] = key_shuffle[4575];
    assign key_original[1671] = key_shuffle[8129];
    assign key_original[1670] = key_shuffle[1500];
    assign key_original[1669] = key_shuffle[2813];
    assign key_original[1668] = key_shuffle[5985];
    assign key_original[1667] = key_shuffle[1033];
    assign key_original[1666] = key_shuffle[6086];
    assign key_original[1665] = key_shuffle[595];
    assign key_original[1664] = key_shuffle[5089];
    assign key_original[1663] = key_shuffle[2056];
    assign key_original[1662] = key_shuffle[1453];
    assign key_original[1661] = key_shuffle[8165];
    assign key_original[1660] = key_shuffle[4475];
    assign key_original[1659] = key_shuffle[76];
    assign key_original[1658] = key_shuffle[6264];
    assign key_original[1657] = key_shuffle[1718];
    assign key_original[1656] = key_shuffle[6719];
    assign key_original[1655] = key_shuffle[7371];
    assign key_original[1654] = key_shuffle[3858];
    assign key_original[1653] = key_shuffle[4334];
    assign key_original[1652] = key_shuffle[5624];
    assign key_original[1651] = key_shuffle[6279];
    assign key_original[1650] = key_shuffle[6492];
    assign key_original[1649] = key_shuffle[5972];
    assign key_original[1648] = key_shuffle[7504];
    assign key_original[1647] = key_shuffle[3782];
    assign key_original[1646] = key_shuffle[7096];
    assign key_original[1645] = key_shuffle[677];
    assign key_original[1644] = key_shuffle[27];
    assign key_original[1643] = key_shuffle[3529];
    assign key_original[1642] = key_shuffle[5594];
    assign key_original[1641] = key_shuffle[6515];
    assign key_original[1640] = key_shuffle[5009];
    assign key_original[1639] = key_shuffle[1025];
    assign key_original[1638] = key_shuffle[7180];
    assign key_original[1637] = key_shuffle[210];
    assign key_original[1636] = key_shuffle[7813];
    assign key_original[1635] = key_shuffle[365];
    assign key_original[1634] = key_shuffle[4325];
    assign key_original[1633] = key_shuffle[7040];
    assign key_original[1632] = key_shuffle[1234];
    assign key_original[1631] = key_shuffle[7165];
    assign key_original[1630] = key_shuffle[7234];
    assign key_original[1629] = key_shuffle[7207];
    assign key_original[1628] = key_shuffle[4332];
    assign key_original[1627] = key_shuffle[713];
    assign key_original[1626] = key_shuffle[5613];
    assign key_original[1625] = key_shuffle[385];
    assign key_original[1624] = key_shuffle[7960];
    assign key_original[1623] = key_shuffle[6579];
    assign key_original[1622] = key_shuffle[2561];
    assign key_original[1621] = key_shuffle[6028];
    assign key_original[1620] = key_shuffle[6924];
    assign key_original[1619] = key_shuffle[6588];
    assign key_original[1618] = key_shuffle[5747];
    assign key_original[1617] = key_shuffle[6484];
    assign key_original[1616] = key_shuffle[3957];
    assign key_original[1615] = key_shuffle[1125];
    assign key_original[1614] = key_shuffle[2713];
    assign key_original[1613] = key_shuffle[351];
    assign key_original[1612] = key_shuffle[6996];
    assign key_original[1611] = key_shuffle[4712];
    assign key_original[1610] = key_shuffle[4692];
    assign key_original[1609] = key_shuffle[3470];
    assign key_original[1608] = key_shuffle[3990];
    assign key_original[1607] = key_shuffle[6316];
    assign key_original[1606] = key_shuffle[1249];
    assign key_original[1605] = key_shuffle[2874];
    assign key_original[1604] = key_shuffle[4493];
    assign key_original[1603] = key_shuffle[5682];
    assign key_original[1602] = key_shuffle[447];
    assign key_original[1601] = key_shuffle[2003];
    assign key_original[1600] = key_shuffle[4893];
    assign key_original[1599] = key_shuffle[5967];
    assign key_original[1598] = key_shuffle[2];
    assign key_original[1597] = key_shuffle[1180];
    assign key_original[1596] = key_shuffle[8085];
    assign key_original[1595] = key_shuffle[670];
    assign key_original[1594] = key_shuffle[3901];
    assign key_original[1593] = key_shuffle[1212];
    assign key_original[1592] = key_shuffle[5360];
    assign key_original[1591] = key_shuffle[4472];
    assign key_original[1590] = key_shuffle[573];
    assign key_original[1589] = key_shuffle[2167];
    assign key_original[1588] = key_shuffle[2042];
    assign key_original[1587] = key_shuffle[4147];
    assign key_original[1586] = key_shuffle[2394];
    assign key_original[1585] = key_shuffle[8122];
    assign key_original[1584] = key_shuffle[2427];
    assign key_original[1583] = key_shuffle[6939];
    assign key_original[1582] = key_shuffle[314];
    assign key_original[1581] = key_shuffle[6464];
    assign key_original[1580] = key_shuffle[8172];
    assign key_original[1579] = key_shuffle[3910];
    assign key_original[1578] = key_shuffle[5402];
    assign key_original[1577] = key_shuffle[6741];
    assign key_original[1576] = key_shuffle[7853];
    assign key_original[1575] = key_shuffle[3840];
    assign key_original[1574] = key_shuffle[4103];
    assign key_original[1573] = key_shuffle[1555];
    assign key_original[1572] = key_shuffle[2718];
    assign key_original[1571] = key_shuffle[7460];
    assign key_original[1570] = key_shuffle[3337];
    assign key_original[1569] = key_shuffle[5450];
    assign key_original[1568] = key_shuffle[7189];
    assign key_original[1567] = key_shuffle[6250];
    assign key_original[1566] = key_shuffle[629];
    assign key_original[1565] = key_shuffle[2537];
    assign key_original[1564] = key_shuffle[693];
    assign key_original[1563] = key_shuffle[3920];
    assign key_original[1562] = key_shuffle[7262];
    assign key_original[1561] = key_shuffle[545];
    assign key_original[1560] = key_shuffle[876];
    assign key_original[1559] = key_shuffle[1960];
    assign key_original[1558] = key_shuffle[6062];
    assign key_original[1557] = key_shuffle[4599];
    assign key_original[1556] = key_shuffle[2138];
    assign key_original[1555] = key_shuffle[6723];
    assign key_original[1554] = key_shuffle[4559];
    assign key_original[1553] = key_shuffle[7715];
    assign key_original[1552] = key_shuffle[1801];
    assign key_original[1551] = key_shuffle[2065];
    assign key_original[1550] = key_shuffle[3941];
    assign key_original[1549] = key_shuffle[6311];
    assign key_original[1548] = key_shuffle[5742];
    assign key_original[1547] = key_shuffle[2209];
    assign key_original[1546] = key_shuffle[4109];
    assign key_original[1545] = key_shuffle[1638];
    assign key_original[1544] = key_shuffle[8184];
    assign key_original[1543] = key_shuffle[6727];
    assign key_original[1542] = key_shuffle[1845];
    assign key_original[1541] = key_shuffle[241];
    assign key_original[1540] = key_shuffle[5138];
    assign key_original[1539] = key_shuffle[8037];
    assign key_original[1538] = key_shuffle[3165];
    assign key_original[1537] = key_shuffle[2805];
    assign key_original[1536] = key_shuffle[7595];
    assign key_original[1535] = key_shuffle[868];
    assign key_original[1534] = key_shuffle[6137];
    assign key_original[1533] = key_shuffle[19];
    assign key_original[1532] = key_shuffle[731];
    assign key_original[1531] = key_shuffle[2071];
    assign key_original[1530] = key_shuffle[1114];
    assign key_original[1529] = key_shuffle[926];
    assign key_original[1528] = key_shuffle[5665];
    assign key_original[1527] = key_shuffle[7638];
    assign key_original[1526] = key_shuffle[1425];
    assign key_original[1525] = key_shuffle[1369];
    assign key_original[1524] = key_shuffle[617];
    assign key_original[1523] = key_shuffle[1600];
    assign key_original[1522] = key_shuffle[73];
    assign key_original[1521] = key_shuffle[7147];
    assign key_original[1520] = key_shuffle[1573];
    assign key_original[1519] = key_shuffle[2973];
    assign key_original[1518] = key_shuffle[5429];
    assign key_original[1517] = key_shuffle[7131];
    assign key_original[1516] = key_shuffle[4686];
    assign key_original[1515] = key_shuffle[7968];
    assign key_original[1514] = key_shuffle[1178];
    assign key_original[1513] = key_shuffle[5897];
    assign key_original[1512] = key_shuffle[5449];
    assign key_original[1511] = key_shuffle[4999];
    assign key_original[1510] = key_shuffle[4055];
    assign key_original[1509] = key_shuffle[6613];
    assign key_original[1508] = key_shuffle[5533];
    assign key_original[1507] = key_shuffle[2062];
    assign key_original[1506] = key_shuffle[6215];
    assign key_original[1505] = key_shuffle[3841];
    assign key_original[1504] = key_shuffle[1368];
    assign key_original[1503] = key_shuffle[409];
    assign key_original[1502] = key_shuffle[5739];
    assign key_original[1501] = key_shuffle[3515];
    assign key_original[1500] = key_shuffle[3104];
    assign key_original[1499] = key_shuffle[2150];
    assign key_original[1498] = key_shuffle[5016];
    assign key_original[1497] = key_shuffle[4];
    assign key_original[1496] = key_shuffle[3549];
    assign key_original[1495] = key_shuffle[4937];
    assign key_original[1494] = key_shuffle[5425];
    assign key_original[1493] = key_shuffle[451];
    assign key_original[1492] = key_shuffle[449];
    assign key_original[1491] = key_shuffle[2357];
    assign key_original[1490] = key_shuffle[5061];
    assign key_original[1489] = key_shuffle[4911];
    assign key_original[1488] = key_shuffle[3183];
    assign key_original[1487] = key_shuffle[7486];
    assign key_original[1486] = key_shuffle[3252];
    assign key_original[1485] = key_shuffle[4084];
    assign key_original[1484] = key_shuffle[4414];
    assign key_original[1483] = key_shuffle[6666];
    assign key_original[1482] = key_shuffle[2141];
    assign key_original[1481] = key_shuffle[7405];
    assign key_original[1480] = key_shuffle[923];
    assign key_original[1479] = key_shuffle[4909];
    assign key_original[1478] = key_shuffle[2407];
    assign key_original[1477] = key_shuffle[6350];
    assign key_original[1476] = key_shuffle[2276];
    assign key_original[1475] = key_shuffle[3987];
    assign key_original[1474] = key_shuffle[3350];
    assign key_original[1473] = key_shuffle[6926];
    assign key_original[1472] = key_shuffle[2885];
    assign key_original[1471] = key_shuffle[1429];
    assign key_original[1470] = key_shuffle[7018];
    assign key_original[1469] = key_shuffle[1014];
    assign key_original[1468] = key_shuffle[5459];
    assign key_original[1467] = key_shuffle[4022];
    assign key_original[1466] = key_shuffle[6814];
    assign key_original[1465] = key_shuffle[1021];
    assign key_original[1464] = key_shuffle[6540];
    assign key_original[1463] = key_shuffle[6781];
    assign key_original[1462] = key_shuffle[7686];
    assign key_original[1461] = key_shuffle[5574];
    assign key_original[1460] = key_shuffle[105];
    assign key_original[1459] = key_shuffle[579];
    assign key_original[1458] = key_shuffle[5908];
    assign key_original[1457] = key_shuffle[5164];
    assign key_original[1456] = key_shuffle[8062];
    assign key_original[1455] = key_shuffle[4955];
    assign key_original[1454] = key_shuffle[6957];
    assign key_original[1453] = key_shuffle[3624];
    assign key_original[1452] = key_shuffle[6005];
    assign key_original[1451] = key_shuffle[2708];
    assign key_original[1450] = key_shuffle[248];
    assign key_original[1449] = key_shuffle[7505];
    assign key_original[1448] = key_shuffle[5346];
    assign key_original[1447] = key_shuffle[5046];
    assign key_original[1446] = key_shuffle[5230];
    assign key_original[1445] = key_shuffle[3399];
    assign key_original[1444] = key_shuffle[3712];
    assign key_original[1443] = key_shuffle[1793];
    assign key_original[1442] = key_shuffle[892];
    assign key_original[1441] = key_shuffle[6868];
    assign key_original[1440] = key_shuffle[3940];
    assign key_original[1439] = key_shuffle[2852];
    assign key_original[1438] = key_shuffle[3625];
    assign key_original[1437] = key_shuffle[3060];
    assign key_original[1436] = key_shuffle[3706];
    assign key_original[1435] = key_shuffle[522];
    assign key_original[1434] = key_shuffle[3604];
    assign key_original[1433] = key_shuffle[3974];
    assign key_original[1432] = key_shuffle[66];
    assign key_original[1431] = key_shuffle[8130];
    assign key_original[1430] = key_shuffle[485];
    assign key_original[1429] = key_shuffle[2909];
    assign key_original[1428] = key_shuffle[202];
    assign key_original[1427] = key_shuffle[4457];
    assign key_original[1426] = key_shuffle[822];
    assign key_original[1425] = key_shuffle[1026];
    assign key_original[1424] = key_shuffle[4337];
    assign key_original[1423] = key_shuffle[2338];
    assign key_original[1422] = key_shuffle[7358];
    assign key_original[1421] = key_shuffle[2865];
    assign key_original[1420] = key_shuffle[1049];
    assign key_original[1419] = key_shuffle[6456];
    assign key_original[1418] = key_shuffle[4584];
    assign key_original[1417] = key_shuffle[4892];
    assign key_original[1416] = key_shuffle[4754];
    assign key_original[1415] = key_shuffle[1451];
    assign key_original[1414] = key_shuffle[7397];
    assign key_original[1413] = key_shuffle[6341];
    assign key_original[1412] = key_shuffle[7141];
    assign key_original[1411] = key_shuffle[2451];
    assign key_original[1410] = key_shuffle[7160];
    assign key_original[1409] = key_shuffle[4293];
    assign key_original[1408] = key_shuffle[3143];
    assign key_original[1407] = key_shuffle[4417];
    assign key_original[1406] = key_shuffle[5752];
    assign key_original[1405] = key_shuffle[1998];
    assign key_original[1404] = key_shuffle[297];
    assign key_original[1403] = key_shuffle[3518];
    assign key_original[1402] = key_shuffle[5465];
    assign key_original[1401] = key_shuffle[5540];
    assign key_original[1400] = key_shuffle[5262];
    assign key_original[1399] = key_shuffle[3370];
    assign key_original[1398] = key_shuffle[6345];
    assign key_original[1397] = key_shuffle[6168];
    assign key_original[1396] = key_shuffle[5782];
    assign key_original[1395] = key_shuffle[57];
    assign key_original[1394] = key_shuffle[3434];
    assign key_original[1393] = key_shuffle[2358];
    assign key_original[1392] = key_shuffle[3816];
    assign key_original[1391] = key_shuffle[1091];
    assign key_original[1390] = key_shuffle[4258];
    assign key_original[1389] = key_shuffle[6692];
    assign key_original[1388] = key_shuffle[5015];
    assign key_original[1387] = key_shuffle[6805];
    assign key_original[1386] = key_shuffle[1350];
    assign key_original[1385] = key_shuffle[4661];
    assign key_original[1384] = key_shuffle[535];
    assign key_original[1383] = key_shuffle[6658];
    assign key_original[1382] = key_shuffle[3167];
    assign key_original[1381] = key_shuffle[5675];
    assign key_original[1380] = key_shuffle[1593];
    assign key_original[1379] = key_shuffle[8133];
    assign key_original[1378] = key_shuffle[5636];
    assign key_original[1377] = key_shuffle[2081];
    assign key_original[1376] = key_shuffle[2344];
    assign key_original[1375] = key_shuffle[7692];
    assign key_original[1374] = key_shuffle[6161];
    assign key_original[1373] = key_shuffle[2773];
    assign key_original[1372] = key_shuffle[6980];
    assign key_original[1371] = key_shuffle[5404];
    assign key_original[1370] = key_shuffle[171];
    assign key_original[1369] = key_shuffle[5826];
    assign key_original[1368] = key_shuffle[5559];
    assign key_original[1367] = key_shuffle[1300];
    assign key_original[1366] = key_shuffle[2514];
    assign key_original[1365] = key_shuffle[6632];
    assign key_original[1364] = key_shuffle[2268];
    assign key_original[1363] = key_shuffle[96];
    assign key_original[1362] = key_shuffle[1649];
    assign key_original[1361] = key_shuffle[2785];
    assign key_original[1360] = key_shuffle[2911];
    assign key_original[1359] = key_shuffle[4344];
    assign key_original[1358] = key_shuffle[368];
    assign key_original[1357] = key_shuffle[1008];
    assign key_original[1356] = key_shuffle[3209];
    assign key_original[1355] = key_shuffle[4825];
    assign key_original[1354] = key_shuffle[4331];
    assign key_original[1353] = key_shuffle[4901];
    assign key_original[1352] = key_shuffle[2461];
    assign key_original[1351] = key_shuffle[705];
    assign key_original[1350] = key_shuffle[2779];
    assign key_original[1349] = key_shuffle[7436];
    assign key_original[1348] = key_shuffle[5471];
    assign key_original[1347] = key_shuffle[3233];
    assign key_original[1346] = key_shuffle[223];
    assign key_original[1345] = key_shuffle[1525];
    assign key_original[1344] = key_shuffle[6116];
    assign key_original[1343] = key_shuffle[6144];
    assign key_original[1342] = key_shuffle[6587];
    assign key_original[1341] = key_shuffle[5397];
    assign key_original[1340] = key_shuffle[7317];
    assign key_original[1339] = key_shuffle[6002];
    assign key_original[1338] = key_shuffle[947];
    assign key_original[1337] = key_shuffle[558];
    assign key_original[1336] = key_shuffle[7193];
    assign key_original[1335] = key_shuffle[6882];
    assign key_original[1334] = key_shuffle[2413];
    assign key_original[1333] = key_shuffle[7870];
    assign key_original[1332] = key_shuffle[5161];
    assign key_original[1331] = key_shuffle[2006];
    assign key_original[1330] = key_shuffle[1677];
    assign key_original[1329] = key_shuffle[7396];
    assign key_original[1328] = key_shuffle[219];
    assign key_original[1327] = key_shuffle[5096];
    assign key_original[1326] = key_shuffle[5505];
    assign key_original[1325] = key_shuffle[185];
    assign key_original[1324] = key_shuffle[7175];
    assign key_original[1323] = key_shuffle[3128];
    assign key_original[1322] = key_shuffle[7824];
    assign key_original[1321] = key_shuffle[3340];
    assign key_original[1320] = key_shuffle[8154];
    assign key_original[1319] = key_shuffle[2360];
    assign key_original[1318] = key_shuffle[8087];
    assign key_original[1317] = key_shuffle[5699];
    assign key_original[1316] = key_shuffle[8071];
    assign key_original[1315] = key_shuffle[7971];
    assign key_original[1314] = key_shuffle[7801];
    assign key_original[1313] = key_shuffle[6174];
    assign key_original[1312] = key_shuffle[5767];
    assign key_original[1311] = key_shuffle[5311];
    assign key_original[1310] = key_shuffle[495];
    assign key_original[1309] = key_shuffle[1557];
    assign key_original[1308] = key_shuffle[3905];
    assign key_original[1307] = key_shuffle[2797];
    assign key_original[1306] = key_shuffle[1292];
    assign key_original[1305] = key_shuffle[3759];
    assign key_original[1304] = key_shuffle[1806];
    assign key_original[1303] = key_shuffle[2674];
    assign key_original[1302] = key_shuffle[588];
    assign key_original[1301] = key_shuffle[7446];
    assign key_original[1300] = key_shuffle[5032];
    assign key_original[1299] = key_shuffle[1496];
    assign key_original[1298] = key_shuffle[1046];
    assign key_original[1297] = key_shuffle[1539];
    assign key_original[1296] = key_shuffle[4320];
    assign key_original[1295] = key_shuffle[2692];
    assign key_original[1294] = key_shuffle[805];
    assign key_original[1293] = key_shuffle[6020];
    assign key_original[1292] = key_shuffle[7297];
    assign key_original[1291] = key_shuffle[6889];
    assign key_original[1290] = key_shuffle[7173];
    assign key_original[1289] = key_shuffle[98];
    assign key_original[1288] = key_shuffle[4544];
    assign key_original[1287] = key_shuffle[3074];
    assign key_original[1286] = key_shuffle[3285];
    assign key_original[1285] = key_shuffle[4391];
    assign key_original[1284] = key_shuffle[5149];
    assign key_original[1283] = key_shuffle[3559];
    assign key_original[1282] = key_shuffle[762];
    assign key_original[1281] = key_shuffle[4890];
    assign key_original[1280] = key_shuffle[1423];
    assign key_original[1279] = key_shuffle[597];
    assign key_original[1278] = key_shuffle[8090];
    assign key_original[1277] = key_shuffle[2947];
    assign key_original[1276] = key_shuffle[823];
    assign key_original[1275] = key_shuffle[181];
    assign key_original[1274] = key_shuffle[878];
    assign key_original[1273] = key_shuffle[3222];
    assign key_original[1272] = key_shuffle[6214];
    assign key_original[1271] = key_shuffle[6787];
    assign key_original[1270] = key_shuffle[2435];
    assign key_original[1269] = key_shuffle[1515];
    assign key_original[1268] = key_shuffle[561];
    assign key_original[1267] = key_shuffle[5889];
    assign key_original[1266] = key_shuffle[4972];
    assign key_original[1265] = key_shuffle[4036];
    assign key_original[1264] = key_shuffle[4633];
    assign key_original[1263] = key_shuffle[2440];
    assign key_original[1262] = key_shuffle[2272];
    assign key_original[1261] = key_shuffle[1280];
    assign key_original[1260] = key_shuffle[827];
    assign key_original[1259] = key_shuffle[1126];
    assign key_original[1258] = key_shuffle[6582];
    assign key_original[1257] = key_shuffle[6033];
    assign key_original[1256] = key_shuffle[7322];
    assign key_original[1255] = key_shuffle[7351];
    assign key_original[1254] = key_shuffle[2551];
    assign key_original[1253] = key_shuffle[4287];
    assign key_original[1252] = key_shuffle[749];
    assign key_original[1251] = key_shuffle[2182];
    assign key_original[1250] = key_shuffle[2719];
    assign key_original[1249] = key_shuffle[2920];
    assign key_original[1248] = key_shuffle[1064];
    assign key_original[1247] = key_shuffle[6353];
    assign key_original[1246] = key_shuffle[3306];
    assign key_original[1245] = key_shuffle[2439];
    assign key_original[1244] = key_shuffle[6700];
    assign key_original[1243] = key_shuffle[4718];
    assign key_original[1242] = key_shuffle[5911];
    assign key_original[1241] = key_shuffle[4595];
    assign key_original[1240] = key_shuffle[3373];
    assign key_original[1239] = key_shuffle[4447];
    assign key_original[1238] = key_shuffle[1371];
    assign key_original[1237] = key_shuffle[20];
    assign key_original[1236] = key_shuffle[3457];
    assign key_original[1235] = key_shuffle[5913];
    assign key_original[1234] = key_shuffle[4555];
    assign key_original[1233] = key_shuffle[5426];
    assign key_original[1232] = key_shuffle[440];
    assign key_original[1231] = key_shuffle[5464];
    assign key_original[1230] = key_shuffle[3194];
    assign key_original[1229] = key_shuffle[4087];
    assign key_original[1228] = key_shuffle[8131];
    assign key_original[1227] = key_shuffle[4698];
    assign key_original[1226] = key_shuffle[4190];
    assign key_original[1225] = key_shuffle[3793];
    assign key_original[1224] = key_shuffle[3689];
    assign key_original[1223] = key_shuffle[6625];
    assign key_original[1222] = key_shuffle[5609];
    assign key_original[1221] = key_shuffle[1383];
    assign key_original[1220] = key_shuffle[4639];
    assign key_original[1219] = key_shuffle[2218];
    assign key_original[1218] = key_shuffle[1459];
    assign key_original[1217] = key_shuffle[1774];
    assign key_original[1216] = key_shuffle[6848];
    assign key_original[1215] = key_shuffle[698];
    assign key_original[1214] = key_shuffle[6057];
    assign key_original[1213] = key_shuffle[1382];
    assign key_original[1212] = key_shuffle[460];
    assign key_original[1211] = key_shuffle[3749];
    assign key_original[1210] = key_shuffle[8086];
    assign key_original[1209] = key_shuffle[7300];
    assign key_original[1208] = key_shuffle[7948];
    assign key_original[1207] = key_shuffle[6241];
    assign key_original[1206] = key_shuffle[2539];
    assign key_original[1205] = key_shuffle[6115];
    assign key_original[1204] = key_shuffle[4214];
    assign key_original[1203] = key_shuffle[3385];
    assign key_original[1202] = key_shuffle[857];
    assign key_original[1201] = key_shuffle[8020];
    assign key_original[1200] = key_shuffle[3734];
    assign key_original[1199] = key_shuffle[5127];
    assign key_original[1198] = key_shuffle[1614];
    assign key_original[1197] = key_shuffle[4183];
    assign key_original[1196] = key_shuffle[4257];
    assign key_original[1195] = key_shuffle[6498];
    assign key_original[1194] = key_shuffle[645];
    assign key_original[1193] = key_shuffle[551];
    assign key_original[1192] = key_shuffle[5191];
    assign key_original[1191] = key_shuffle[5165];
    assign key_original[1190] = key_shuffle[5258];
    assign key_original[1189] = key_shuffle[5359];
    assign key_original[1188] = key_shuffle[1154];
    assign key_original[1187] = key_shuffle[6544];
    assign key_original[1186] = key_shuffle[1331];
    assign key_original[1185] = key_shuffle[5833];
    assign key_original[1184] = key_shuffle[3973];
    assign key_original[1183] = key_shuffle[5135];
    assign key_original[1182] = key_shuffle[1595];
    assign key_original[1181] = key_shuffle[1812];
    assign key_original[1180] = key_shuffle[5483];
    assign key_original[1179] = key_shuffle[3438];
    assign key_original[1178] = key_shuffle[6773];
    assign key_original[1177] = key_shuffle[5381];
    assign key_original[1176] = key_shuffle[6758];
    assign key_original[1175] = key_shuffle[5303];
    assign key_original[1174] = key_shuffle[5700];
    assign key_original[1173] = key_shuffle[3444];
    assign key_original[1172] = key_shuffle[2682];
    assign key_original[1171] = key_shuffle[2125];
    assign key_original[1170] = key_shuffle[3287];
    assign key_original[1169] = key_shuffle[5677];
    assign key_original[1168] = key_shuffle[7064];
    assign key_original[1167] = key_shuffle[8142];
    assign key_original[1166] = key_shuffle[1147];
    assign key_original[1165] = key_shuffle[6881];
    assign key_original[1164] = key_shuffle[5620];
    assign key_original[1163] = key_shuffle[6517];
    assign key_original[1162] = key_shuffle[5881];
    assign key_original[1161] = key_shuffle[88];
    assign key_original[1160] = key_shuffle[2233];
    assign key_original[1159] = key_shuffle[7417];
    assign key_original[1158] = key_shuffle[3207];
    assign key_original[1157] = key_shuffle[7875];
    assign key_original[1156] = key_shuffle[4570];
    assign key_original[1155] = key_shuffle[2907];
    assign key_original[1154] = key_shuffle[6626];
    assign key_original[1153] = key_shuffle[6334];
    assign key_original[1152] = key_shuffle[676];
    assign key_original[1151] = key_shuffle[1495];
    assign key_original[1150] = key_shuffle[4360];
    assign key_original[1149] = key_shuffle[2541];
    assign key_original[1148] = key_shuffle[1524];
    assign key_original[1147] = key_shuffle[6995];
    assign key_original[1146] = key_shuffle[1824];
    assign key_original[1145] = key_shuffle[7836];
    assign key_original[1144] = key_shuffle[3929];
    assign key_original[1143] = key_shuffle[7600];
    assign key_original[1142] = key_shuffle[1951];
    assign key_original[1141] = key_shuffle[5673];
    assign key_original[1140] = key_shuffle[7266];
    assign key_original[1139] = key_shuffle[7273];
    assign key_original[1138] = key_shuffle[1517];
    assign key_original[1137] = key_shuffle[6536];
    assign key_original[1136] = key_shuffle[2825];
    assign key_original[1135] = key_shuffle[7626];
    assign key_original[1134] = key_shuffle[345];
    assign key_original[1133] = key_shuffle[4756];
    assign key_original[1132] = key_shuffle[306];
    assign key_original[1131] = key_shuffle[3288];
    assign key_original[1130] = key_shuffle[3154];
    assign key_original[1129] = key_shuffle[1431];
    assign key_original[1128] = key_shuffle[1494];
    assign key_original[1127] = key_shuffle[4424];
    assign key_original[1126] = key_shuffle[7336];
    assign key_original[1125] = key_shuffle[7622];
    assign key_original[1124] = key_shuffle[7541];
    assign key_original[1123] = key_shuffle[6771];
    assign key_original[1122] = key_shuffle[6474];
    assign key_original[1121] = key_shuffle[7657];
    assign key_original[1120] = key_shuffle[114];
    assign key_original[1119] = key_shuffle[8136];
    assign key_original[1118] = key_shuffle[3907];
    assign key_original[1117] = key_shuffle[941];
    assign key_original[1116] = key_shuffle[785];
    assign key_original[1115] = key_shuffle[7606];
    assign key_original[1114] = key_shuffle[3994];
    assign key_original[1113] = key_shuffle[6813];
    assign key_original[1112] = key_shuffle[2099];
    assign key_original[1111] = key_shuffle[7445];
    assign key_original[1110] = key_shuffle[2817];
    assign key_original[1109] = key_shuffle[6550];
    assign key_original[1108] = key_shuffle[2023];
    assign key_original[1107] = key_shuffle[2002];
    assign key_original[1106] = key_shuffle[5734];
    assign key_original[1105] = key_shuffle[3717];
    assign key_original[1104] = key_shuffle[6876];
    assign key_original[1103] = key_shuffle[3486];
    assign key_original[1102] = key_shuffle[6034];
    assign key_original[1101] = key_shuffle[6208];
    assign key_original[1100] = key_shuffle[4211];
    assign key_original[1099] = key_shuffle[1137];
    assign key_original[1098] = key_shuffle[2203];
    assign key_original[1097] = key_shuffle[3641];
    assign key_original[1096] = key_shuffle[1645];
    assign key_original[1095] = key_shuffle[2273];
    assign key_original[1094] = key_shuffle[1190];
    assign key_original[1093] = key_shuffle[6179];
    assign key_original[1092] = key_shuffle[56];
    assign key_original[1091] = key_shuffle[968];
    assign key_original[1090] = key_shuffle[608];
    assign key_original[1089] = key_shuffle[3334];
    assign key_original[1088] = key_shuffle[307];
    assign key_original[1087] = key_shuffle[6731];
    assign key_original[1086] = key_shuffle[1699];
    assign key_original[1085] = key_shuffle[7103];
    assign key_original[1084] = key_shuffle[811];
    assign key_original[1083] = key_shuffle[6642];
    assign key_original[1082] = key_shuffle[5770];
    assign key_original[1081] = key_shuffle[2853];
    assign key_original[1080] = key_shuffle[7529];
    assign key_original[1079] = key_shuffle[2041];
    assign key_original[1078] = key_shuffle[7972];
    assign key_original[1077] = key_shuffle[641];
    assign key_original[1076] = key_shuffle[1311];
    assign key_original[1075] = key_shuffle[7623];
    assign key_original[1074] = key_shuffle[4437];
    assign key_original[1073] = key_shuffle[1417];
    assign key_original[1072] = key_shuffle[3672];
    assign key_original[1071] = key_shuffle[549];
    assign key_original[1070] = key_shuffle[2396];
    assign key_original[1069] = key_shuffle[7897];
    assign key_original[1068] = key_shuffle[7557];
    assign key_original[1067] = key_shuffle[740];
    assign key_original[1066] = key_shuffle[5308];
    assign key_original[1065] = key_shuffle[72];
    assign key_original[1064] = key_shuffle[4159];
    assign key_original[1063] = key_shuffle[6159];
    assign key_original[1062] = key_shuffle[309];
    assign key_original[1061] = key_shuffle[1173];
    assign key_original[1060] = key_shuffle[1612];
    assign key_original[1059] = key_shuffle[6981];
    assign key_original[1058] = key_shuffle[7602];
    assign key_original[1057] = key_shuffle[4834];
    assign key_original[1056] = key_shuffle[1585];
    assign key_original[1055] = key_shuffle[5909];
    assign key_original[1054] = key_shuffle[7292];
    assign key_original[1053] = key_shuffle[921];
    assign key_original[1052] = key_shuffle[3397];
    assign key_original[1051] = key_shuffle[2673];
    assign key_original[1050] = key_shuffle[6987];
    assign key_original[1049] = key_shuffle[5413];
    assign key_original[1048] = key_shuffle[5649];
    assign key_original[1047] = key_shuffle[4425];
    assign key_original[1046] = key_shuffle[2492];
    assign key_original[1045] = key_shuffle[186];
    assign key_original[1044] = key_shuffle[1825];
    assign key_original[1043] = key_shuffle[1219];
    assign key_original[1042] = key_shuffle[1281];
    assign key_original[1041] = key_shuffle[6669];
    assign key_original[1040] = key_shuffle[1732];
    assign key_original[1039] = key_shuffle[7673];
    assign key_original[1038] = key_shuffle[674];
    assign key_original[1037] = key_shuffle[3521];
    assign key_original[1036] = key_shuffle[1606];
    assign key_original[1035] = key_shuffle[3058];
    assign key_original[1034] = key_shuffle[4523];
    assign key_original[1033] = key_shuffle[1908];
    assign key_original[1032] = key_shuffle[5731];
    assign key_original[1031] = key_shuffle[5436];
    assign key_original[1030] = key_shuffle[1118];
    assign key_original[1029] = key_shuffle[6156];
    assign key_original[1028] = key_shuffle[2925];
    assign key_original[1027] = key_shuffle[381];
    assign key_original[1026] = key_shuffle[7143];
    assign key_original[1025] = key_shuffle[1839];
    assign key_original[1024] = key_shuffle[7572];
    assign key_original[1023] = key_shuffle[1017];
    assign key_original[1022] = key_shuffle[4614];
    assign key_original[1021] = key_shuffle[6003];
    assign key_original[1020] = key_shuffle[251];
    assign key_original[1019] = key_shuffle[6902];
    assign key_original[1018] = key_shuffle[4900];
    assign key_original[1017] = key_shuffle[7896];
    assign key_original[1016] = key_shuffle[7803];
    assign key_original[1015] = key_shuffle[7343];
    assign key_original[1014] = key_shuffle[4647];
    assign key_original[1013] = key_shuffle[7681];
    assign key_original[1012] = key_shuffle[7823];
    assign key_original[1011] = key_shuffle[2311];
    assign key_original[1010] = key_shuffle[4156];
    assign key_original[1009] = key_shuffle[425];
    assign key_original[1008] = key_shuffle[2212];
    assign key_original[1007] = key_shuffle[4566];
    assign key_original[1006] = key_shuffle[4586];
    assign key_original[1005] = key_shuffle[5433];
    assign key_original[1004] = key_shuffle[4792];
    assign key_original[1003] = key_shuffle[2285];
    assign key_original[1002] = key_shuffle[7261];
    assign key_original[1001] = key_shuffle[2742];
    assign key_original[1000] = key_shuffle[2838];
    assign key_original[999] = key_shuffle[5845];
    assign key_original[998] = key_shuffle[5188];
    assign key_original[997] = key_shuffle[5097];
    assign key_original[996] = key_shuffle[8064];
    assign key_original[995] = key_shuffle[7523];
    assign key_original[994] = key_shuffle[7901];
    assign key_original[993] = key_shuffle[3532];
    assign key_original[992] = key_shuffle[5237];
    assign key_original[991] = key_shuffle[2487];
    assign key_original[990] = key_shuffle[298];
    assign key_original[989] = key_shuffle[3912];
    assign key_original[988] = key_shuffle[432];
    assign key_original[987] = key_shuffle[646];
    assign key_original[986] = key_shuffle[5668];
    assign key_original[985] = key_shuffle[6411];
    assign key_original[984] = key_shuffle[8134];
    assign key_original[983] = key_shuffle[7402];
    assign key_original[982] = key_shuffle[7475];
    assign key_original[981] = key_shuffle[543];
    assign key_original[980] = key_shuffle[5332];
    assign key_original[979] = key_shuffle[4120];
    assign key_original[978] = key_shuffle[6825];
    assign key_original[977] = key_shuffle[5374];
    assign key_original[976] = key_shuffle[4831];
    assign key_original[975] = key_shuffle[1742];
    assign key_original[974] = key_shuffle[5380];
    assign key_original[973] = key_shuffle[6918];
    assign key_original[972] = key_shuffle[4784];
    assign key_original[971] = key_shuffle[1725];
    assign key_original[970] = key_shuffle[1295];
    assign key_original[969] = key_shuffle[4564];
    assign key_original[968] = key_shuffle[801];
    assign key_original[967] = key_shuffle[6932];
    assign key_original[966] = key_shuffle[5705];
    assign key_original[965] = key_shuffle[4198];
    assign key_original[964] = key_shuffle[2807];
    assign key_original[963] = key_shuffle[667];
    assign key_original[962] = key_shuffle[4311];
    assign key_original[961] = key_shuffle[5882];
    assign key_original[960] = key_shuffle[424];
    assign key_original[959] = key_shuffle[1379];
    assign key_original[958] = key_shuffle[5761];
    assign key_original[957] = key_shuffle[5940];
    assign key_original[956] = key_shuffle[1140];
    assign key_original[955] = key_shuffle[5802];
    assign key_original[954] = key_shuffle[2074];
    assign key_original[953] = key_shuffle[7226];
    assign key_original[952] = key_shuffle[4627];
    assign key_original[951] = key_shuffle[1558];
    assign key_original[950] = key_shuffle[7170];
    assign key_original[949] = key_shuffle[1222];
    assign key_original[948] = key_shuffle[3786];
    assign key_original[947] = key_shuffle[7166];
    assign key_original[946] = key_shuffle[4206];
    assign key_original[945] = key_shuffle[592];
    assign key_original[944] = key_shuffle[139];
    assign key_original[943] = key_shuffle[5725];
    assign key_original[942] = key_shuffle[812];
    assign key_original[941] = key_shuffle[1225];
    assign key_original[940] = key_shuffle[3344];
    assign key_original[939] = key_shuffle[8027];
    assign key_original[938] = key_shuffle[5905];
    assign key_original[937] = key_shuffle[5275];
    assign key_original[936] = key_shuffle[6195];
    assign key_original[935] = key_shuffle[3915];
    assign key_original[934] = key_shuffle[4889];
    assign key_original[933] = key_shuffle[7962];
    assign key_original[932] = key_shuffle[3900];
    assign key_original[931] = key_shuffle[2446];
    assign key_original[930] = key_shuffle[1692];
    assign key_original[929] = key_shuffle[1727];
    assign key_original[928] = key_shuffle[5888];
    assign key_original[927] = key_shuffle[696];
    assign key_original[926] = key_shuffle[6392];
    assign key_original[925] = key_shuffle[4050];
    assign key_original[924] = key_shuffle[457];
    assign key_original[923] = key_shuffle[3576];
    assign key_original[922] = key_shuffle[4781];
    assign key_original[921] = key_shuffle[4220];
    assign key_original[920] = key_shuffle[3366];
    assign key_original[919] = key_shuffle[6489];
    assign key_original[918] = key_shuffle[7357];
    assign key_original[917] = key_shuffle[1018];
    assign key_original[916] = key_shuffle[416];
    assign key_original[915] = key_shuffle[5547];
    assign key_original[914] = key_shuffle[2130];
    assign key_original[913] = key_shuffle[7146];
    assign key_original[912] = key_shuffle[5110];
    assign key_original[911] = key_shuffle[998];
    assign key_original[910] = key_shuffle[1213];
    assign key_original[909] = key_shuffle[7366];
    assign key_original[908] = key_shuffle[3417];
    assign key_original[907] = key_shuffle[5176];
    assign key_original[906] = key_shuffle[2493];
    assign key_original[905] = key_shuffle[235];
    assign key_original[904] = key_shuffle[7565];
    assign key_original[903] = key_shuffle[2980];
    assign key_original[902] = key_shuffle[4942];
    assign key_original[901] = key_shuffle[4603];
    assign key_original[900] = key_shuffle[2555];
    assign key_original[899] = key_shuffle[258];
    assign key_original[898] = key_shuffle[6499];
    assign key_original[897] = key_shuffle[2022];
    assign key_original[896] = key_shuffle[2686];
    assign key_original[895] = key_shuffle[4796];
    assign key_original[894] = key_shuffle[1589];
    assign key_original[893] = key_shuffle[5104];
    assign key_original[892] = key_shuffle[2077];
    assign key_original[891] = key_shuffle[1165];
    assign key_original[890] = key_shuffle[6344];
    assign key_original[889] = key_shuffle[62];
    assign key_original[888] = key_shuffle[1401];
    assign key_original[887] = key_shuffle[807];
    assign key_original[886] = key_shuffle[3155];
    assign key_original[885] = key_shuffle[2417];
    assign key_original[884] = key_shuffle[6574];
    assign key_original[883] = key_shuffle[7301];
    assign key_original[882] = key_shuffle[4797];
    assign key_original[881] = key_shuffle[51];
    assign key_original[880] = key_shuffle[4019];
    assign key_original[879] = key_shuffle[3355];
    assign key_original[878] = key_shuffle[8187];
    assign key_original[877] = key_shuffle[302];
    assign key_original[876] = key_shuffle[7025];
    assign key_original[875] = key_shuffle[771];
    assign key_original[874] = key_shuffle[7002];
    assign key_original[873] = key_shuffle[3797];
    assign key_original[872] = key_shuffle[6473];
    assign key_original[871] = key_shuffle[2712];
    assign key_original[870] = key_shuffle[3919];
    assign key_original[869] = key_shuffle[8153];
    assign key_original[868] = key_shuffle[6035];
    assign key_original[867] = key_shuffle[418];
    assign key_original[866] = key_shuffle[3335];
    assign key_original[865] = key_shuffle[5589];
    assign key_original[864] = key_shuffle[1983];
    assign key_original[863] = key_shuffle[4759];
    assign key_original[862] = key_shuffle[2012];
    assign key_original[861] = key_shuffle[6313];
    assign key_original[860] = key_shuffle[1623];
    assign key_original[859] = key_shuffle[6716];
    assign key_original[858] = key_shuffle[1358];
    assign key_original[857] = key_shuffle[1167];
    assign key_original[856] = key_shuffle[5553];
    assign key_original[855] = key_shuffle[7593];
    assign key_original[854] = key_shuffle[3217];
    assign key_original[853] = key_shuffle[7133];
    assign key_original[852] = key_shuffle[6670];
    assign key_original[851] = key_shuffle[4454];
    assign key_original[850] = key_shuffle[7211];
    assign key_original[849] = key_shuffle[8186];
    assign key_original[848] = key_shuffle[2049];
    assign key_original[847] = key_shuffle[4520];
    assign key_original[846] = key_shuffle[5345];
    assign key_original[845] = key_shuffle[971];
    assign key_original[844] = key_shuffle[2271];
    assign key_original[843] = key_shuffle[8023];
    assign key_original[842] = key_shuffle[1858];
    assign key_original[841] = key_shuffle[7735];
    assign key_original[840] = key_shuffle[854];
    assign key_original[839] = key_shuffle[7876];
    assign key_original[838] = key_shuffle[3032];
    assign key_original[837] = key_shuffle[1899];
    assign key_original[836] = key_shuffle[3918];
    assign key_original[835] = key_shuffle[4151];
    assign key_original[834] = key_shuffle[4587];
    assign key_original[833] = key_shuffle[4277];
    assign key_original[832] = key_shuffle[1688];
    assign key_original[831] = key_shuffle[1363];
    assign key_original[830] = key_shuffle[7974];
    assign key_original[829] = key_shuffle[3849];
    assign key_original[828] = key_shuffle[2899];
    assign key_original[827] = key_shuffle[6067];
    assign key_original[826] = key_shuffle[4021];
    assign key_original[825] = key_shuffle[4116];
    assign key_original[824] = key_shuffle[2126];
    assign key_original[823] = key_shuffle[789];
    assign key_original[822] = key_shuffle[2111];
    assign key_original[821] = key_shuffle[2464];
    assign key_original[820] = key_shuffle[5143];
    assign key_original[819] = key_shuffle[3286];
    assign key_original[818] = key_shuffle[5645];
    assign key_original[817] = key_shuffle[3455];
    assign key_original[816] = key_shuffle[2731];
    assign key_original[815] = key_shuffle[4172];
    assign key_original[814] = key_shuffle[8137];
    assign key_original[813] = key_shuffle[1741];
    assign key_original[812] = key_shuffle[5638];
    assign key_original[811] = key_shuffle[7831];
    assign key_original[810] = key_shuffle[4928];
    assign key_original[809] = key_shuffle[7553];
    assign key_original[808] = key_shuffle[3550];
    assign key_original[807] = key_shuffle[3179];
    assign key_original[806] = key_shuffle[4229];
    assign key_original[805] = key_shuffle[5883];
    assign key_original[804] = key_shuffle[4958];
    assign key_original[803] = key_shuffle[902];
    assign key_original[802] = key_shuffle[1993];
    assign key_original[801] = key_shuffle[6896];
    assign key_original[800] = key_shuffle[7094];
    assign key_original[799] = key_shuffle[7755];
    assign key_original[798] = key_shuffle[688];
    assign key_original[797] = key_shuffle[7710];
    assign key_original[796] = key_shuffle[1491];
    assign key_original[795] = key_shuffle[1526];
    assign key_original[794] = key_shuffle[6355];
    assign key_original[793] = key_shuffle[7409];
    assign key_original[792] = key_shuffle[2050];
    assign key_original[791] = key_shuffle[330];
    assign key_original[790] = key_shuffle[6095];
    assign key_original[789] = key_shuffle[3139];
    assign key_original[788] = key_shuffle[2101];
    assign key_original[787] = key_shuffle[85];
    assign key_original[786] = key_shuffle[7142];
    assign key_original[785] = key_shuffle[6739];
    assign key_original[784] = key_shuffle[3828];
    assign key_original[783] = key_shuffle[2476];
    assign key_original[782] = key_shuffle[395];
    assign key_original[781] = key_shuffle[2132];
    assign key_original[780] = key_shuffle[8115];
    assign key_original[779] = key_shuffle[3251];
    assign key_original[778] = key_shuffle[2337];
    assign key_original[777] = key_shuffle[3788];
    assign key_original[776] = key_shuffle[3160];
    assign key_original[775] = key_shuffle[1995];
    assign key_original[774] = key_shuffle[6122];
    assign key_original[773] = key_shuffle[5339];
    assign key_original[772] = key_shuffle[2053];
    assign key_original[771] = key_shuffle[6906];
    assign key_original[770] = key_shuffle[1990];
    assign key_original[769] = key_shuffle[1115];
    assign key_original[768] = key_shuffle[2191];
    assign key_original[767] = key_shuffle[4908];
    assign key_original[766] = key_shuffle[5510];
    assign key_original[765] = key_shuffle[4905];
    assign key_original[764] = key_shuffle[5995];
    assign key_original[763] = key_shuffle[4435];
    assign key_original[762] = key_shuffle[4826];
    assign key_original[761] = key_shuffle[2059];
    assign key_original[760] = key_shuffle[1963];
    assign key_original[759] = key_shuffle[2110];
    assign key_original[758] = key_shuffle[150];
    assign key_original[757] = key_shuffle[555];
    assign key_original[756] = key_shuffle[6864];
    assign key_original[755] = key_shuffle[3906];
    assign key_original[754] = key_shuffle[3193];
    assign key_original[753] = key_shuffle[2609];
    assign key_original[752] = key_shuffle[2113];
    assign key_original[751] = key_shuffle[624];
    assign key_original[750] = key_shuffle[2955];
    assign key_original[749] = key_shuffle[7576];
    assign key_original[748] = key_shuffle[5331];
    assign key_original[747] = key_shuffle[2129];
    assign key_original[746] = key_shuffle[5861];
    assign key_original[745] = key_shuffle[5541];
    assign key_original[744] = key_shuffle[7411];
    assign key_original[743] = key_shuffle[4551];
    assign key_original[742] = key_shuffle[6472];
    assign key_original[741] = key_shuffle[7346];
    assign key_original[740] = key_shuffle[927];
    assign key_original[739] = key_shuffle[6628];
    assign key_original[738] = key_shuffle[5565];
    assign key_original[737] = key_shuffle[8088];
    assign key_original[736] = key_shuffle[4481];
    assign key_original[735] = key_shuffle[4939];
    assign key_original[734] = key_shuffle[2240];
    assign key_original[733] = key_shuffle[7152];
    assign key_original[732] = key_shuffle[7369];
    assign key_original[731] = key_shuffle[4176];
    assign key_original[730] = key_shuffle[858];
    assign key_original[729] = key_shuffle[3720];
    assign key_original[728] = key_shuffle[4256];
    assign key_original[727] = key_shuffle[7124];
    assign key_original[726] = key_shuffle[2324];
    assign key_original[725] = key_shuffle[7167];
    assign key_original[724] = key_shuffle[3618];
    assign key_original[723] = key_shuffle[1866];
    assign key_original[722] = key_shuffle[1669];
    assign key_original[721] = key_shuffle[3181];
    assign key_original[720] = key_shuffle[2675];
    assign key_original[719] = key_shuffle[1723];
    assign key_original[718] = key_shuffle[612];
    assign key_original[717] = key_shuffle[5003];
    assign key_original[716] = key_shuffle[1586];
    assign key_original[715] = key_shuffle[4582];
    assign key_original[714] = key_shuffle[4767];
    assign key_original[713] = key_shuffle[6610];
    assign key_original[712] = key_shuffle[8073];
    assign key_original[711] = key_shuffle[313];
    assign key_original[710] = key_shuffle[3493];
    assign key_original[709] = key_shuffle[8024];
    assign key_original[708] = key_shuffle[4716];
    assign key_original[707] = key_shuffle[4588];
    assign key_original[706] = key_shuffle[2669];
    assign key_original[705] = key_shuffle[1504];
    assign key_original[704] = key_shuffle[3320];
    assign key_original[703] = key_shuffle[6450];
    assign key_original[702] = key_shuffle[3188];
    assign key_original[701] = key_shuffle[3378];
    assign key_original[700] = key_shuffle[7691];
    assign key_original[699] = key_shuffle[67];
    assign key_original[698] = key_shuffle[4572];
    assign key_original[697] = key_shuffle[4996];
    assign key_original[696] = key_shuffle[6835];
    assign key_original[695] = key_shuffle[7527];
    assign key_original[694] = key_shuffle[249];
    assign key_original[693] = key_shuffle[6007];
    assign key_original[692] = key_shuffle[108];
    assign key_original[691] = key_shuffle[3784];
    assign key_original[690] = key_shuffle[3092];
    assign key_original[689] = key_shuffle[1454];
    assign key_original[688] = key_shuffle[5103];
    assign key_original[687] = key_shuffle[865];
    assign key_original[686] = key_shuffle[6196];
    assign key_original[685] = key_shuffle[2275];
    assign key_original[684] = key_shuffle[1072];
    assign key_original[683] = key_shuffle[2607];
    assign key_original[682] = key_shuffle[104];
    assign key_original[681] = key_shuffle[5685];
    assign key_original[680] = key_shuffle[2703];
    assign key_original[679] = key_shuffle[1894];
    assign key_original[678] = key_shuffle[7482];
    assign key_original[677] = key_shuffle[2162];
    assign key_original[676] = key_shuffle[4702];
    assign key_original[675] = key_shuffle[5693];
    assign key_original[674] = key_shuffle[4506];
    assign key_original[673] = key_shuffle[7634];
    assign key_original[672] = key_shuffle[4944];
    assign key_original[671] = key_shuffle[7121];
    assign key_original[670] = key_shuffle[6754];
    assign key_original[669] = key_shuffle[301];
    assign key_original[668] = key_shuffle[2291];
    assign key_original[667] = key_shuffle[1928];
    assign key_original[666] = key_shuffle[5282];
    assign key_original[665] = key_shuffle[4253];
    assign key_original[664] = key_shuffle[3351];
    assign key_original[663] = key_shuffle[5643];
    assign key_original[662] = key_shuffle[236];
    assign key_original[661] = key_shuffle[4141];
    assign key_original[660] = key_shuffle[1925];
    assign key_original[659] = key_shuffle[1922];
    assign key_original[658] = key_shuffle[1550];
    assign key_original[657] = key_shuffle[1119];
    assign key_original[656] = key_shuffle[6999];
    assign key_original[655] = key_shuffle[152];
    assign key_original[654] = key_shuffle[3197];
    assign key_original[653] = key_shuffle[1706];
    assign key_original[652] = key_shuffle[3191];
    assign key_original[651] = key_shuffle[2072];
    assign key_original[650] = key_shuffle[7182];
    assign key_original[649] = key_shuffle[6520];
    assign key_original[648] = key_shuffle[2371];
    assign key_original[647] = key_shuffle[5492];
    assign key_original[646] = key_shuffle[8093];
    assign key_original[645] = key_shuffle[402];
    assign key_original[644] = key_shuffle[3667];
    assign key_original[643] = key_shuffle[7291];
    assign key_original[642] = key_shuffle[1261];
    assign key_original[641] = key_shuffle[3673];
    assign key_original[640] = key_shuffle[1888];
    assign key_original[639] = key_shuffle[6445];
    assign key_original[638] = key_shuffle[572];
    assign key_original[637] = key_shuffle[1215];
    assign key_original[636] = key_shuffle[2981];
    assign key_original[635] = key_shuffle[4177];
    assign key_original[634] = key_shuffle[3614];
    assign key_original[633] = key_shuffle[3086];
    assign key_original[632] = key_shuffle[6463];
    assign key_original[631] = key_shuffle[5177];
    assign key_original[630] = key_shuffle[1544];
    assign key_original[629] = key_shuffle[4399];
    assign key_original[628] = key_shuffle[4817];
    assign key_original[627] = key_shuffle[2032];
    assign key_original[626] = key_shuffle[178];
    assign key_original[625] = key_shuffle[3296];
    assign key_original[624] = key_shuffle[3897];
    assign key_original[623] = key_shuffle[5587];
    assign key_original[622] = key_shuffle[864];
    assign key_original[621] = key_shuffle[835];
    assign key_original[620] = key_shuffle[7992];
    assign key_original[619] = key_shuffle[958];
    assign key_original[618] = key_shuffle[623];
    assign key_original[617] = key_shuffle[506];
    assign key_original[616] = key_shuffle[6618];
    assign key_original[615] = key_shuffle[841];
    assign key_original[614] = key_shuffle[4690];
    assign key_original[613] = key_shuffle[3503];
    assign key_original[612] = key_shuffle[7407];
    assign key_original[611] = key_shuffle[5997];
    assign key_original[610] = key_shuffle[4850];
    assign key_original[609] = key_shuffle[149];
    assign key_original[608] = key_shuffle[593];
    assign key_original[607] = key_shuffle[1411];
    assign key_original[606] = key_shuffle[6629];
    assign key_original[605] = key_shuffle[2013];
    assign key_original[604] = key_shuffle[2530];
    assign key_original[603] = key_shuffle[63];
    assign key_original[602] = key_shuffle[2466];
    assign key_original[601] = key_shuffle[3605];
    assign key_original[600] = key_shuffle[7574];
    assign key_original[599] = key_shuffle[3998];
    assign key_original[598] = key_shuffle[5328];
    assign key_original[597] = key_shuffle[6711];
    assign key_original[596] = key_shuffle[6875];
    assign key_original[595] = key_shuffle[5156];
    assign key_original[594] = key_shuffle[3441];
    assign key_original[593] = key_shuffle[949];
    assign key_original[592] = key_shuffle[5812];
    assign key_original[591] = key_shuffle[4025];
    assign key_original[590] = key_shuffle[6160];
    assign key_original[589] = key_shuffle[7422];
    assign key_original[588] = key_shuffle[5158];
    assign key_original[587] = key_shuffle[93];
    assign key_original[586] = key_shuffle[5651];
    assign key_original[585] = key_shuffle[466];
    assign key_original[584] = key_shuffle[5715];
    assign key_original[583] = key_shuffle[3298];
    assign key_original[582] = key_shuffle[6139];
    assign key_original[581] = key_shuffle[5460];
    assign key_original[580] = key_shuffle[2327];
    assign key_original[579] = key_shuffle[1245];
    assign key_original[578] = key_shuffle[6269];
    assign key_original[577] = key_shuffle[4795];
    assign key_original[576] = key_shuffle[1354];
    assign key_original[575] = key_shuffle[6127];
    assign key_original[574] = key_shuffle[4473];
    assign key_original[573] = key_shuffle[2892];
    assign key_original[572] = key_shuffle[6880];
    assign key_original[571] = key_shuffle[340];
    assign key_original[570] = key_shuffle[5961];
    assign key_original[569] = key_shuffle[734];
    assign key_original[568] = key_shuffle[3156];
    assign key_original[567] = key_shuffle[836];
    assign key_original[566] = key_shuffle[3108];
    assign key_original[565] = key_shuffle[7398];
    assign key_original[564] = key_shuffle[5674];
    assign key_original[563] = key_shuffle[172];
    assign key_original[562] = key_shuffle[5593];
    assign key_original[561] = key_shuffle[4057];
    assign key_original[560] = key_shuffle[1789];
    assign key_original[559] = key_shuffle[5671];
    assign key_original[558] = key_shuffle[3416];
    assign key_original[557] = key_shuffle[7621];
    assign key_original[556] = key_shuffle[2747];
    assign key_original[555] = key_shuffle[2502];
    assign key_original[554] = key_shuffle[3813];
    assign key_original[553] = key_shuffle[4123];
    assign key_original[552] = key_shuffle[400];
    assign key_original[551] = key_shuffle[2567];
    assign key_original[550] = key_shuffle[1150];
    assign key_original[549] = key_shuffle[4298];
    assign key_original[548] = key_shuffle[7325];
    assign key_original[547] = key_shuffle[2559];
    assign key_original[546] = key_shuffle[6190];
    assign key_original[545] = key_shuffle[2355];
    assign key_original[544] = key_shuffle[7042];
    assign key_original[543] = key_shuffle[4010];
    assign key_original[542] = key_shuffle[3305];
    assign key_original[541] = key_shuffle[1492];
    assign key_original[540] = key_shuffle[1498];
    assign key_original[539] = key_shuffle[3668];
    assign key_original[538] = key_shuffle[5270];
    assign key_original[537] = key_shuffle[3362];
    assign key_original[536] = key_shuffle[7179];
    assign key_original[535] = key_shuffle[2603];
    assign key_original[534] = key_shuffle[1989];
    assign key_original[533] = key_shuffle[7660];
    assign key_original[532] = key_shuffle[2670];
    assign key_original[531] = key_shuffle[6584];
    assign key_original[530] = key_shuffle[6266];
    assign key_original[529] = key_shuffle[1207];
    assign key_original[528] = key_shuffle[2334];
    assign key_original[527] = key_shuffle[4170];
    assign key_original[526] = key_shuffle[8135];
    assign key_original[525] = key_shuffle[6091];
    assign key_original[524] = key_shuffle[1887];
    assign key_original[523] = key_shuffle[4415];
    assign key_original[522] = key_shuffle[5720];
    assign key_original[521] = key_shuffle[113];
    assign key_original[520] = key_shuffle[7232];
    assign key_original[519] = key_shuffle[1136];
    assign key_original[518] = key_shuffle[6583];
    assign key_original[517] = key_shuffle[3684];
    assign key_original[516] = key_shuffle[6227];
    assign key_original[515] = key_shuffle[3501];
    assign key_original[514] = key_shuffle[1107];
    assign key_original[513] = key_shuffle[4442];
    assign key_original[512] = key_shuffle[3293];
    assign key_original[511] = key_shuffle[1608];
    assign key_original[510] = key_shuffle[6972];
    assign key_original[509] = key_shuffle[3246];
    assign key_original[508] = key_shuffle[4730];
    assign key_original[507] = key_shuffle[2608];
    assign key_original[506] = key_shuffle[5386];
    assign key_original[505] = key_shuffle[1944];
    assign key_original[504] = key_shuffle[1932];
    assign key_original[503] = key_shuffle[4122];
    assign key_original[502] = key_shuffle[7985];
    assign key_original[501] = key_shuffle[5867];
    assign key_original[500] = key_shuffle[6274];
    assign key_original[499] = key_shuffle[5874];
    assign key_original[498] = key_shuffle[1821];
    assign key_original[497] = key_shuffle[4226];
    assign key_original[496] = key_shuffle[1452];
    assign key_original[495] = key_shuffle[1755];
    assign key_original[494] = key_shuffle[1621];
    assign key_original[493] = key_shuffle[1591];
    assign key_original[492] = key_shuffle[7473];
    assign key_original[491] = key_shuffle[183];
    assign key_original[490] = key_shuffle[5515];
    assign key_original[489] = key_shuffle[7868];
    assign key_original[488] = key_shuffle[4413];
    assign key_original[487] = key_shuffle[6408];
    assign key_original[486] = key_shuffle[754];
    assign key_original[485] = key_shuffle[7811];
    assign key_original[484] = key_shuffle[1315];
    assign key_original[483] = key_shuffle[7923];
    assign key_original[482] = key_shuffle[4461];
    assign key_original[481] = key_shuffle[905];
    assign key_original[480] = key_shuffle[1923];
    assign key_original[479] = key_shuffle[954];
    assign key_original[478] = key_shuffle[1179];
    assign key_original[477] = key_shuffle[7187];
    assign key_original[476] = key_shuffle[5748];
    assign key_original[475] = key_shuffle[2465];
    assign key_original[474] = key_shuffle[4460];
    assign key_original[473] = key_shuffle[4090];
    assign key_original[472] = key_shuffle[3872];
    assign key_original[471] = key_shuffle[5033];
    assign key_original[470] = key_shuffle[3279];
    assign key_original[469] = key_shuffle[7395];
    assign key_original[468] = key_shuffle[3471];
    assign key_original[467] = key_shuffle[4101];
    assign key_original[466] = key_shuffle[278];
    assign key_original[465] = key_shuffle[222];
    assign key_original[464] = key_shuffle[2657];
    assign key_original[463] = key_shuffle[3925];
    assign key_original[462] = key_shuffle[4394];
    assign key_original[461] = key_shuffle[7852];
    assign key_original[460] = key_shuffle[6529];
    assign key_original[459] = key_shuffle[1533];
    assign key_original[458] = key_shuffle[601];
    assign key_original[457] = key_shuffle[6085];
    assign key_original[456] = key_shuffle[7288];
    assign key_original[455] = key_shuffle[3376];
    assign key_original[454] = key_shuffle[7507];
    assign key_original[453] = key_shuffle[8005];
    assign key_original[452] = key_shuffle[1768];
    assign key_original[451] = key_shuffle[2858];
    assign key_original[450] = key_shuffle[8052];
    assign key_original[449] = key_shuffle[5052];
    assign key_original[448] = key_shuffle[3753];
    assign key_original[447] = key_shuffle[167];
    assign key_original[446] = key_shuffle[2136];
    assign key_original[445] = key_shuffle[3324];
    assign key_original[444] = key_shuffle[4887];
    assign key_original[443] = key_shuffle[2565];
    assign key_original[442] = key_shuffle[7698];
    assign key_original[441] = key_shuffle[6760];
    assign key_original[440] = key_shuffle[7684];
    assign key_original[439] = key_shuffle[862];
    assign key_original[438] = key_shuffle[4636];
    assign key_original[437] = key_shuffle[195];
    assign key_original[436] = key_shuffle[3675];
    assign key_original[435] = key_shuffle[3939];
    assign key_original[434] = key_shuffle[2710];
    assign key_original[433] = key_shuffle[2905];
    assign key_original[432] = key_shuffle[2821];
    assign key_original[431] = key_shuffle[3853];
    assign key_original[430] = key_shuffle[2769];
    assign key_original[429] = key_shuffle[5984];
    assign key_original[428] = key_shuffle[7869];
    assign key_original[427] = key_shuffle[1009];
    assign key_original[426] = key_shuffle[2749];
    assign key_original[425] = key_shuffle[609];
    assign key_original[424] = key_shuffle[3175];
    assign key_original[423] = key_shuffle[1276];
    assign key_original[422] = key_shuffle[7864];
    assign key_original[421] = key_shuffle[6125];
    assign key_original[420] = key_shuffle[111];
    assign key_original[419] = key_shuffle[3875];
    assign key_original[418] = key_shuffle[7194];
    assign key_original[417] = key_shuffle[1301];
    assign key_original[416] = key_shuffle[6979];
    assign key_original[415] = key_shuffle[4770];
    assign key_original[414] = key_shuffle[3890];
    assign key_original[413] = key_shuffle[2880];
    assign key_original[412] = key_shuffle[8049];
    assign key_original[411] = key_shuffle[3770];
    assign key_original[410] = key_shuffle[2794];
    assign key_original[409] = key_shuffle[5575];
    assign key_original[408] = key_shuffle[4524];
    assign key_original[407] = key_shuffle[7725];
    assign key_original[406] = key_shuffle[5486];
    assign key_original[405] = key_shuffle[2962];
    assign key_original[404] = key_shuffle[4094];
    assign key_original[403] = key_shuffle[619];
    assign key_original[402] = key_shuffle[95];
    assign key_original[401] = key_shuffle[6560];
    assign key_original[400] = key_shuffle[2726];
    assign key_original[399] = key_shuffle[5115];
    assign key_original[398] = key_shuffle[5523];
    assign key_original[397] = key_shuffle[7704];
    assign key_original[396] = key_shuffle[1715];
    assign key_original[395] = key_shuffle[6737];
    assign key_original[394] = key_shuffle[7385];
    assign key_original[393] = key_shuffle[7466];
    assign key_original[392] = key_shuffle[6808];
    assign key_original[391] = key_shuffle[6884];
    assign key_original[390] = key_shuffle[6207];
    assign key_original[389] = key_shuffle[4228];
    assign key_original[388] = key_shuffle[5820];
    assign key_original[387] = key_shuffle[5169];
    assign key_original[386] = key_shuffle[6024];
    assign key_original[385] = key_shuffle[82];
    assign key_original[384] = key_shuffle[5903];
    assign key_original[383] = key_shuffle[4538];
    assign key_original[382] = key_shuffle[5468];
    assign key_original[381] = key_shuffle[8067];
    assign key_original[380] = key_shuffle[4201];
    assign key_original[379] = key_shuffle[1877];
    assign key_original[378] = key_shuffle[1782];
    assign key_original[377] = key_shuffle[2227];
    assign key_original[376] = key_shuffle[5773];
    assign key_original[375] = key_shuffle[2035];
    assign key_original[374] = key_shuffle[41];
    assign key_original[373] = key_shuffle[3884];
    assign key_original[372] = key_shuffle[4745];
    assign key_original[371] = key_shuffle[1584];
    assign key_original[370] = key_shuffle[5774];
    assign key_original[369] = key_shuffle[3682];
    assign key_original[368] = key_shuffle[6487];
    assign key_original[367] = key_shuffle[3547];
    assign key_original[366] = key_shuffle[7248];
    assign key_original[365] = key_shuffle[5930];
    assign key_original[364] = key_shuffle[4724];
    assign key_original[363] = key_shuffle[3001];
    assign key_original[362] = key_shuffle[7904];
    assign key_original[361] = key_shuffle[3028];
    assign key_original[360] = key_shuffle[1353];
    assign key_original[359] = key_shuffle[738];
    assign key_original[358] = key_shuffle[1603];
    assign key_original[357] = key_shuffle[453];
    assign key_original[356] = key_shuffle[564];
    assign key_original[355] = key_shuffle[2245];
    assign key_original[354] = key_shuffle[7871];
    assign key_original[353] = key_shuffle[3100];
    assign key_original[352] = key_shuffle[4175];
    assign key_original[351] = key_shuffle[4691];
    assign key_original[350] = key_shuffle[6083];
    assign key_original[349] = key_shuffle[169];
    assign key_original[348] = key_shuffle[5444];
    assign key_original[347] = key_shuffle[4707];
    assign key_original[346] = key_shuffle[7975];
    assign key_original[345] = key_shuffle[5178];
    assign key_original[344] = key_shuffle[7082];
    assign key_original[343] = key_shuffle[4670];
    assign key_original[342] = key_shuffle[4780];
    assign key_original[341] = key_shuffle[7675];
    assign key_original[340] = key_shuffle[651];
    assign key_original[339] = key_shuffle[7521];
    assign key_original[338] = key_shuffle[2063];
    assign key_original[337] = key_shuffle[7027];
    assign key_original[336] = key_shuffle[5746];
    assign key_original[335] = key_shuffle[4933];
    assign key_original[334] = key_shuffle[6585];
    assign key_original[333] = key_shuffle[3484];
    assign key_original[332] = key_shuffle[6998];
    assign key_original[331] = key_shuffle[6636];
    assign key_original[330] = key_shuffle[6436];
    assign key_original[329] = key_shuffle[1783];
    assign key_original[328] = key_shuffle[7547];
    assign key_original[327] = key_shuffle[1911];
    assign key_original[326] = key_shuffle[2527];
    assign key_original[325] = key_shuffle[4338];
    assign key_original[324] = key_shuffle[2632];
    assign key_original[323] = key_shuffle[5470];
    assign key_original[322] = key_shuffle[1132];
    assign key_original[321] = key_shuffle[7073];
    assign key_original[320] = key_shuffle[2257];
    assign key_original[319] = key_shuffle[3114];
    assign key_original[318] = key_shuffle[5482];
    assign key_original[317] = key_shuffle[3826];
    assign key_original[316] = key_shuffle[174];
    assign key_original[315] = key_shuffle[631];
    assign key_original[314] = key_shuffle[6494];
    assign key_original[313] = key_shuffle[5676];
    assign key_original[312] = key_shuffle[2140];
    assign key_original[311] = key_shuffle[3377];
    assign key_original[310] = key_shuffle[4187];
    assign key_original[309] = key_shuffle[3119];
    assign key_original[308] = key_shuffle[3023];
    assign key_original[307] = key_shuffle[2549];
    assign key_original[306] = key_shuffle[2277];
    assign key_original[305] = key_shuffle[2288];
    assign key_original[304] = key_shuffle[658];
    assign key_original[303] = key_shuffle[4728];
    assign key_original[302] = key_shuffle[5088];
    assign key_original[301] = key_shuffle[7635];
    assign key_original[300] = key_shuffle[6405];
    assign key_original[299] = key_shuffle[7826];
    assign key_original[298] = key_shuffle[1881];
    assign key_original[297] = key_shuffle[7646];
    assign key_original[296] = key_shuffle[7973];
    assign key_original[295] = key_shuffle[5252];
    assign key_original[294] = key_shuffle[4153];
    assign key_original[293] = key_shuffle[1113];
    assign key_original[292] = key_shuffle[6521];
    assign key_original[291] = key_shuffle[7344];
    assign key_original[290] = key_shuffle[4593];
    assign key_original[289] = key_shuffle[1659];
    assign key_original[288] = key_shuffle[8162];
    assign key_original[287] = key_shuffle[1055];
    assign key_original[286] = key_shuffle[7873];
    assign key_original[285] = key_shuffle[491];
    assign key_original[284] = key_shuffle[840];
    assign key_original[283] = key_shuffle[3888];
    assign key_original[282] = key_shuffle[2307];
    assign key_original[281] = key_shuffle[7902];
    assign key_original[280] = key_shuffle[3661];
    assign key_original[279] = key_shuffle[2765];
    assign key_original[278] = key_shuffle[4567];
    assign key_original[277] = key_shuffle[6129];
    assign key_original[276] = key_shuffle[2993];
    assign key_original[275] = key_shuffle[3403];
    assign key_original[274] = key_shuffle[4312];
    assign key_original[273] = key_shuffle[343];
    assign key_original[272] = key_shuffle[2771];
    assign key_original[271] = key_shuffle[5785];
    assign key_original[270] = key_shuffle[6853];
    assign key_original[269] = key_shuffle[7178];
    assign key_original[268] = key_shuffle[1386];
    assign key_original[267] = key_shuffle[242];
    assign key_original[266] = key_shuffle[7506];
    assign key_original[265] = key_shuffle[5738];
    assign key_original[264] = key_shuffle[3146];
    assign key_original[263] = key_shuffle[5647];
    assign key_original[262] = key_shuffle[5836];
    assign key_original[261] = key_shuffle[218];
    assign key_original[260] = key_shuffle[4818];
    assign key_original[259] = key_shuffle[1419];
    assign key_original[258] = key_shuffle[8032];
    assign key_original[257] = key_shuffle[6885];
    assign key_original[256] = key_shuffle[4852];
    assign key_original[255] = key_shuffle[406];
    assign key_original[254] = key_shuffle[6280];
    assign key_original[253] = key_shuffle[7563];
    assign key_original[252] = key_shuffle[6638];
    assign key_original[251] = key_shuffle[1838];
    assign key_original[250] = key_shuffle[7268];
    assign key_original[249] = key_shuffle[127];
    assign key_original[248] = key_shuffle[2263];
    assign key_original[247] = key_shuffle[1879];
    assign key_original[246] = key_shuffle[335];
    assign key_original[245] = key_shuffle[3835];
    assign key_original[244] = key_shuffle[1474];
    assign key_original[243] = key_shuffle[7849];
    assign key_original[242] = key_shuffle[8177];
    assign key_original[241] = key_shuffle[3459];
    assign key_original[240] = key_shuffle[925];
    assign key_original[239] = key_shuffle[3442];
    assign key_original[238] = key_shuffle[5280];
    assign key_original[237] = key_shuffle[6306];
    assign key_original[236] = key_shuffle[8077];
    assign key_original[235] = key_shuffle[1288];
    assign key_original[234] = key_shuffle[7410];
    assign key_original[233] = key_shuffle[2246];
    assign key_original[232] = key_shuffle[5522];
    assign key_original[231] = key_shuffle[1469];
    assign key_original[230] = key_shuffle[1702];
    assign key_original[229] = key_shuffle[2546];
    assign key_original[228] = key_shuffle[3273];
    assign key_original[227] = key_shuffle[4979];
    assign key_original[226] = key_shuffle[5623];
    assign key_original[225] = key_shuffle[1105];
    assign key_original[224] = key_shuffle[6171];
    assign key_original[223] = key_shuffle[7767];
    assign key_original[222] = key_shuffle[4907];
    assign key_original[221] = key_shuffle[4498];
    assign key_original[220] = key_shuffle[4169];
    assign key_original[219] = key_shuffle[5281];
    assign key_original[218] = key_shuffle[5759];
    assign key_original[217] = key_shuffle[4758];
    assign key_original[216] = key_shuffle[5238];
    assign key_original[215] = key_shuffle[6154];
    assign key_original[214] = key_shuffle[2210];
    assign key_original[213] = key_shuffle[299];
    assign key_original[212] = key_shuffle[5044];
    assign key_original[211] = key_shuffle[4392];
    assign key_original[210] = key_shuffle[919];
    assign key_original[209] = key_shuffle[2028];
    assign key_original[208] = key_shuffle[6495];
    assign key_original[207] = key_shuffle[1422];
    assign key_original[206] = key_shuffle[7746];
    assign key_original[205] = key_shuffle[2998];
    assign key_original[204] = key_shuffle[5163];
    assign key_original[203] = key_shuffle[4964];
    assign key_original[202] = key_shuffle[7403];
    assign key_original[201] = key_shuffle[1704];
    assign key_original[200] = key_shuffle[2626];
    assign key_original[199] = key_shuffle[7881];
    assign key_original[198] = key_shuffle[367];
    assign key_original[197] = key_shuffle[1836];
    assign key_original[196] = key_shuffle[4200];
    assign key_original[195] = key_shuffle[3692];
    assign key_original[194] = key_shuffle[3663];
    assign key_original[193] = key_shuffle[5993];
    assign key_original[192] = key_shuffle[8158];
    assign key_original[191] = key_shuffle[322];
    assign key_original[190] = key_shuffle[4616];
    assign key_original[189] = key_shuffle[481];
    assign key_original[188] = key_shuffle[4056];
    assign key_original[187] = key_shuffle[1689];
    assign key_original[186] = key_shuffle[1316];
    assign key_original[185] = key_shuffle[5198];
    assign key_original[184] = key_shuffle[5914];
    assign key_original[183] = key_shuffle[5606];
    assign key_original[182] = key_shuffle[7821];
    assign key_original[181] = key_shuffle[2701];
    assign key_original[180] = key_shuffle[2634];
    assign key_original[179] = key_shuffle[6282];
    assign key_original[178] = key_shuffle[7014];
    assign key_original[177] = key_shuffle[7947];
    assign key_original[176] = key_shuffle[4932];
    assign key_original[175] = key_shuffle[3328];
    assign key_original[174] = key_shuffle[5255];
    assign key_original[173] = key_shuffle[4791];
    assign key_original[172] = key_shuffle[6372];
    assign key_original[171] = key_shuffle[7356];
    assign key_original[170] = key_shuffle[5692];
    assign key_original[169] = key_shuffle[1643];
    assign key_original[168] = key_shuffle[2877];
    assign key_original[167] = key_shuffle[6175];
    assign key_original[166] = key_shuffle[2621];
    assign key_original[165] = key_shuffle[4925];
    assign key_original[164] = key_shuffle[802];
    assign key_original[163] = key_shuffle[7102];
    assign key_original[162] = key_shuffle[3476];
    assign key_original[161] = key_shuffle[6325];
    assign key_original[160] = key_shuffle[4803];
    assign key_original[159] = key_shuffle[1948];
    assign key_original[158] = key_shuffle[3127];
    assign key_original[157] = key_shuffle[473];
    assign key_original[156] = key_shuffle[7640];
    assign key_original[155] = key_shuffle[2207];
    assign key_original[154] = key_shuffle[5278];
    assign key_original[153] = key_shuffle[4193];
    assign key_original[152] = key_shuffle[5751];
    assign key_original[151] = key_shuffle[7805];
    assign key_original[150] = key_shuffle[8040];
    assign key_original[149] = key_shuffle[2582];
    assign key_original[148] = key_shuffle[7911];
    assign key_original[147] = key_shuffle[1143];
    assign key_original[146] = key_shuffle[965];
    assign key_original[145] = key_shuffle[3043];
    assign key_original[144] = key_shuffle[5251];
    assign key_original[143] = key_shuffle[2937];
    assign key_original[142] = key_shuffle[1152];
    assign key_original[141] = key_shuffle[6539];
    assign key_original[140] = key_shuffle[1720];
    assign key_original[139] = key_shuffle[7361];
    assign key_original[138] = key_shuffle[7799];
    assign key_original[137] = key_shuffle[3943];
    assign key_original[136] = key_shuffle[7855];
    assign key_original[135] = key_shuffle[3313];
    assign key_original[134] = key_shuffle[5557];
    assign key_original[133] = key_shuffle[6414];
    assign key_original[132] = key_shuffle[3634];
    assign key_original[131] = key_shuffle[3769];
    assign key_original[130] = key_shuffle[3019];
    assign key_original[129] = key_shuffle[6049];
    assign key_original[128] = key_shuffle[4967];
    assign key_original[127] = key_shuffle[2406];
    assign key_original[126] = key_shuffle[1760];
    assign key_original[125] = key_shuffle[5023];
    assign key_original[124] = key_shuffle[2721];
    assign key_original[123] = key_shuffle[445];
    assign key_original[122] = key_shuffle[3435];
    assign key_original[121] = key_shuffle[422];
    assign key_original[120] = key_shuffle[315];
    assign key_original[119] = key_shuffle[1442];
    assign key_original[118] = key_shuffle[1096];
    assign key_original[117] = key_shuffle[5101];
    assign key_original[116] = key_shuffle[2055];
    assign key_original[115] = key_shuffle[4003];
    assign key_original[114] = key_shuffle[1788];
    assign key_original[113] = key_shuffle[2823];
    assign key_original[112] = key_shuffle[1362];
    assign key_original[111] = key_shuffle[2971];
    assign key_original[110] = key_shuffle[4263];
    assign key_original[109] = key_shuffle[3781];
    assign key_original[108] = key_shuffle[7932];
    assign key_original[107] = key_shuffle[7037];
    assign key_original[106] = key_shuffle[6103];
    assign key_original[105] = key_shuffle[6772];
    assign key_original[104] = key_shuffle[7671];
    assign key_original[103] = key_shuffle[2664];
    assign key_original[102] = key_shuffle[4063];
    assign key_original[101] = key_shuffle[7987];
    assign key_original[100] = key_shuffle[7424];
    assign key_original[99] = key_shuffle[2420];
    assign key_original[98] = key_shuffle[7499];
    assign key_original[97] = key_shuffle[1334];
    assign key_original[96] = key_shuffle[871];
    assign key_original[95] = key_shuffle[3530];
    assign key_original[94] = key_shuffle[6572];
    assign key_original[93] = key_shuffle[5749];
    assign key_original[92] = key_shuffle[4916];
    assign key_original[91] = key_shuffle[477];
    assign key_original[90] = key_shuffle[344];
    assign key_original[89] = key_shuffle[3047];
    assign key_original[88] = key_shuffle[2562];
    assign key_original[87] = key_shuffle[7748];
    assign key_original[86] = key_shuffle[325];
    assign key_original[85] = key_shuffle[955];
    assign key_original[84] = key_shuffle[5786];
    assign key_original[83] = key_shuffle[6268];
    assign key_original[82] = key_shuffle[7046];
    assign key_original[81] = key_shuffle[1556];
    assign key_original[80] = key_shuffle[3643];
    assign key_original[79] = key_shuffle[2036];
    assign key_original[78] = key_shuffle[7427];
    assign key_original[77] = key_shuffle[5375];
    assign key_original[76] = key_shuffle[2037];
    assign key_original[75] = key_shuffle[672];
    assign key_original[74] = key_shuffle[1694];
    assign key_original[73] = key_shuffle[2881];
    assign key_original[72] = key_shuffle[1841];
    assign key_original[71] = key_shuffle[5393];
    assign key_original[70] = key_shuffle[6821];
    assign key_original[69] = key_shuffle[7625];
    assign key_original[68] = key_shuffle[2158];
    assign key_original[67] = key_shuffle[1996];
    assign key_original[66] = key_shuffle[1882];
    assign key_original[65] = key_shuffle[6229];
    assign key_original[64] = key_shuffle[2419];
    assign key_original[63] = key_shuffle[2982];
    assign key_original[62] = key_shuffle[4291];
    assign key_original[61] = key_shuffle[6479];
    assign key_original[60] = key_shuffle[2016];
    assign key_original[59] = key_shuffle[3846];
    assign key_original[58] = key_shuffle[7525];
    assign key_original[57] = key_shuffle[4534];
    assign key_original[56] = key_shuffle[6132];
    assign key_original[55] = key_shuffle[1283];
    assign key_original[54] = key_shuffle[1785];
    assign key_original[53] = key_shuffle[787];
    assign key_original[52] = key_shuffle[3522];
    assign key_original[51] = key_shuffle[3463];
    assign key_original[50] = key_shuffle[6141];
    assign key_original[49] = key_shuffle[6222];
    assign key_original[48] = key_shuffle[311];
    assign key_original[47] = key_shuffle[3379];
    assign key_original[46] = key_shuffle[3055];
    assign key_original[45] = key_shuffle[7429];
    assign key_original[44] = key_shuffle[4071];
    assign key_original[43] = key_shuffle[1238];
    assign key_original[42] = key_shuffle[461];
    assign key_original[41] = key_shuffle[1461];
    assign key_original[40] = key_shuffle[3574];
    assign key_original[39] = key_shuffle[7782];
    assign key_original[38] = key_shuffle[3636];
    assign key_original[37] = key_shuffle[611];
    assign key_original[36] = key_shuffle[2737];
    assign key_original[35] = key_shuffle[1290];
    assign key_original[34] = key_shuffle[1228];
    assign key_original[33] = key_shuffle[7761];
    assign key_original[32] = key_shuffle[6909];
    assign key_original[31] = key_shuffle[6928];
    assign key_original[30] = key_shuffle[3052];
    assign key_original[29] = key_shuffle[6575];
    assign key_original[28] = key_shuffle[2671];
    assign key_original[27] = key_shuffle[5202];
    assign key_original[26] = key_shuffle[2068];
    assign key_original[25] = key_shuffle[7983];
    assign key_original[24] = key_shuffle[7169];
    assign key_original[23] = key_shuffle[7834];
    assign key_original[22] = key_shuffle[2935];
    assign key_original[21] = key_shuffle[621];
    assign key_original[20] = key_shuffle[2928];
    assign key_original[19] = key_shuffle[1853];
    assign key_original[18] = key_shuffle[1693];
    assign key_original[17] = key_shuffle[3088];
    assign key_original[16] = key_shuffle[1392];
    assign key_original[15] = key_shuffle[5980];
    assign key_original[14] = key_shuffle[4136];
    assign key_original[13] = key_shuffle[4089];
    assign key_original[12] = key_shuffle[7909];
    assign key_original[11] = key_shuffle[5819];
    assign key_original[10] = key_shuffle[590];
    assign key_original[9] = key_shuffle[2428];
    assign key_original[8] = key_shuffle[2760];
    assign key_original[7] = key_shuffle[3494];
    assign key_original[6] = key_shuffle[725];
    assign key_original[5] = key_shuffle[7450];
    assign key_original[4] = key_shuffle[1581];
    assign key_original[3] = key_shuffle[5712];
    assign key_original[2] = key_shuffle[6978];
    assign key_original[1] = key_shuffle[3243];
    assign key_original[0] = key_shuffle[5004];

endmodule