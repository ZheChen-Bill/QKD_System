

//1229 * 36
//36 word length
//32 fraction length


module log2_p_table(
    input [11-1:0] index, //0~2047
    output reg [36-1:0] table_out //36 word length, 32 fraction length
);

    always @(*) begin
        case (index)
            11'd0: table_out = 36'hf4369373b;
            11'd1: table_out = 36'hf438fac0d;
            11'd2: table_out = 36'hf43b61cdd;
            11'd3: table_out = 36'hf43dc89ae;
            11'd4: table_out = 36'hf4402f280;
            11'd5: table_out = 36'hf44295753;
            11'd6: table_out = 36'hf444fb82a;
            11'd7: table_out = 36'hf44761503;
            11'd8: table_out = 36'hf449c6de1;
            11'd9: table_out = 36'hf44c2c2c5;
            11'd10: table_out = 36'hf44e913ae;
            11'd11: table_out = 36'hf450f609e;
            11'd12: table_out = 36'hf4535a995;
            11'd13: table_out = 36'hf455bee95;
            11'd14: table_out = 36'hf45822f9f;
            11'd15: table_out = 36'hf45a86cb2;
            11'd16: table_out = 36'hf45cea5d0;
            11'd17: table_out = 36'hf45f4dafa;
            11'd18: table_out = 36'hf461b0c31;
            11'd19: table_out = 36'hf46413974;
            11'd20: table_out = 36'hf466762c6;
            11'd21: table_out = 36'hf468d8827;
            11'd22: table_out = 36'hf46b3a998;
            11'd23: table_out = 36'hf46d9c71a;
            11'd24: table_out = 36'hf46ffe0ac;
            11'd25: table_out = 36'hf4725f651;
            11'd26: table_out = 36'hf474c080a;
            11'd27: table_out = 36'hf477215d5;
            11'd28: table_out = 36'hf47981fb6;
            11'd29: table_out = 36'hf47be25ac;
            11'd30: table_out = 36'hf47e427b8;
            11'd31: table_out = 36'hf480a25dc;
            11'd32: table_out = 36'hf48302017;
            11'd33: table_out = 36'hf4856166b;
            11'd34: table_out = 36'hf487c08d9;
            11'd35: table_out = 36'hf48a1f760;
            11'd36: table_out = 36'hf48c7e203;
            11'd37: table_out = 36'hf48edc8c2;
            11'd38: table_out = 36'hf4913ab9d;
            11'd39: table_out = 36'hf49398a96;
            11'd40: table_out = 36'hf495f65ad;
            11'd41: table_out = 36'hf49853ce4;
            11'd42: table_out = 36'hf49ab103a;
            11'd43: table_out = 36'hf49d0dfb0;
            11'd44: table_out = 36'hf49f6ab49;
            11'd45: table_out = 36'hf4a1c7303;
            11'd46: table_out = 36'hf4a4236e1;
            11'd47: table_out = 36'hf4a67f6e2;
            11'd48: table_out = 36'hf4a8db308;
            11'd49: table_out = 36'hf4ab36b53;
            11'd50: table_out = 36'hf4ad91fc5;
            11'd51: table_out = 36'hf4afed05d;
            11'd52: table_out = 36'hf4b247d1d;
            11'd53: table_out = 36'hf4b4a2606;
            11'd54: table_out = 36'hf4b6fcb18;
            11'd55: table_out = 36'hf4b956c55;
            11'd56: table_out = 36'hf4bbb09bc;
            11'd57: table_out = 36'hf4be0a34f;
            11'd58: table_out = 36'hf4c06390e;
            11'd59: table_out = 36'hf4c2bcafa;
            11'd60: table_out = 36'hf4c515915;
            11'd61: table_out = 36'hf4c76e35e;
            11'd62: table_out = 36'hf4c9c69d7;
            11'd63: table_out = 36'hf4cc1ec80;
            11'd64: table_out = 36'hf4ce76b5b;
            11'd65: table_out = 36'hf4d0ce667;
            11'd66: table_out = 36'hf4d325da6;
            11'd67: table_out = 36'hf4d57d118;
            11'd68: table_out = 36'hf4d7d40be;
            11'd69: table_out = 36'hf4da2ac9a;
            11'd70: table_out = 36'hf4dc814ab;
            11'd71: table_out = 36'hf4ded78f2;
            11'd72: table_out = 36'hf4e12d971;
            11'd73: table_out = 36'hf4e383628;
            11'd74: table_out = 36'hf4e5d8f18;
            11'd75: table_out = 36'hf4e82e441;
            11'd76: table_out = 36'hf4ea835a5;
            11'd77: table_out = 36'hf4ecd8344;
            11'd78: table_out = 36'hf4ef2cd1e;
            11'd79: table_out = 36'hf4f181335;
            11'd80: table_out = 36'hf4f3d558a;
            11'd81: table_out = 36'hf4f62941c;
            11'd82: table_out = 36'hf4f87ceee;
            11'd83: table_out = 36'hf4fad05ff;
            11'd84: table_out = 36'hf4fd23951;
            11'd85: table_out = 36'hf4ff768e3;
            11'd86: table_out = 36'hf501c94b8;
            11'd87: table_out = 36'hf5041bccf;
            11'd88: table_out = 36'hf5066e12a;
            11'd89: table_out = 36'hf508c01c9;
            11'd90: table_out = 36'hf50b11eac;
            11'd91: table_out = 36'hf50d637d6;
            11'd92: table_out = 36'hf50fb4d46;
            11'd93: table_out = 36'hf51205efd;
            11'd94: table_out = 36'hf51456cfb;
            11'd95: table_out = 36'hf516a7743;
            11'd96: table_out = 36'hf518f7dd4;
            11'd97: table_out = 36'hf51b480af;
            11'd98: table_out = 36'hf51d97fd5;
            11'd99: table_out = 36'hf51fe7b46;
            11'd100: table_out = 36'hf52237304;
            11'd101: table_out = 36'hf5248670f;
            11'd102: table_out = 36'hf526d5768;
            11'd103: table_out = 36'hf52924410;
            11'd104: table_out = 36'hf52b72d06;
            11'd105: table_out = 36'hf52dc124d;
            11'd106: table_out = 36'hf5300f3e5;
            11'd107: table_out = 36'hf5325d1ce;
            11'd108: table_out = 36'hf534aac09;
            11'd109: table_out = 36'hf536f8298;
            11'd110: table_out = 36'hf5394557a;
            11'd111: table_out = 36'hf53b924b1;
            11'd112: table_out = 36'hf53ddf03c;
            11'd113: table_out = 36'hf5402b81e;
            11'd114: table_out = 36'hf54277c57;
            11'd115: table_out = 36'hf544c3ce6;
            11'd116: table_out = 36'hf5470f9ce;
            11'd117: table_out = 36'hf5495b30f;
            11'd118: table_out = 36'hf54ba68a9;
            11'd119: table_out = 36'hf54df1a9e;
            11'd120: table_out = 36'hf5503c8ed;
            11'd121: table_out = 36'hf55287399;
            11'd122: table_out = 36'hf554d1aa1;
            11'd123: table_out = 36'hf5571be06;
            11'd124: table_out = 36'hf55965dc9;
            11'd125: table_out = 36'hf55baf9ea;
            11'd126: table_out = 36'hf55df926b;
            11'd127: table_out = 36'hf5604274c;
            11'd128: table_out = 36'hf5628b88e;
            11'd129: table_out = 36'hf564d4631;
            11'd130: table_out = 36'hf5671d036;
            11'd131: table_out = 36'hf5696569f;
            11'd132: table_out = 36'hf56bad96b;
            11'd133: table_out = 36'hf56df589b;
            11'd134: table_out = 36'hf5703d430;
            11'd135: table_out = 36'hf57284c2c;
            11'd136: table_out = 36'hf574cc08d;
            11'd137: table_out = 36'hf57713156;
            11'd138: table_out = 36'hf57959e87;
            11'd139: table_out = 36'hf57ba0821;
            11'd140: table_out = 36'hf57de6e23;
            11'd141: table_out = 36'hf5802d090;
            11'd142: table_out = 36'hf58272f68;
            11'd143: table_out = 36'hf584b8aab;
            11'd144: table_out = 36'hf586fe25a;
            11'd145: table_out = 36'hf58943676;
            11'd146: table_out = 36'hf58b88700;
            11'd147: table_out = 36'hf58dcd3f8;
            11'd148: table_out = 36'hf59011d5e;
            11'd149: table_out = 36'hf59256335;
            11'd150: table_out = 36'hf5949a57c;
            11'd151: table_out = 36'hf596de434;
            11'd152: table_out = 36'hf59921f5d;
            11'd153: table_out = 36'hf59b656f9;
            11'd154: table_out = 36'hf59da8b09;
            11'd155: table_out = 36'hf59febb8c;
            11'd156: table_out = 36'hf5a22e884;
            11'd157: table_out = 36'hf5a4711f1;
            11'd158: table_out = 36'hf5a6b37d3;
            11'd159: table_out = 36'hf5a8f5a2d;
            11'd160: table_out = 36'hf5ab378fe;
            11'd161: table_out = 36'hf5ad79447;
            11'd162: table_out = 36'hf5afbac08;
            11'd163: table_out = 36'hf5b1fc043;
            11'd164: table_out = 36'hf5b43d0f8;
            11'd165: table_out = 36'hf5b67de28;
            11'd166: table_out = 36'hf5b8be7d3;
            11'd167: table_out = 36'hf5bafedfa;
            11'd168: table_out = 36'hf5bd3f09e;
            11'd169: table_out = 36'hf5bf7efc0;
            11'd170: table_out = 36'hf5c1beb60;
            11'd171: table_out = 36'hf5c3fe37f;
            11'd172: table_out = 36'hf5c63d81d;
            11'd173: table_out = 36'hf5c87c93c;
            11'd174: table_out = 36'hf5cabb6db;
            11'd175: table_out = 36'hf5ccfa0fc;
            11'd176: table_out = 36'hf5cf3879f;
            11'd177: table_out = 36'hf5d176ac6;
            11'd178: table_out = 36'hf5d3b4a70;
            11'd179: table_out = 36'hf5d5f269e;
            11'd180: table_out = 36'hf5d82ff51;
            11'd181: table_out = 36'hf5da6d48a;
            11'd182: table_out = 36'hf5dcaa649;
            11'd183: table_out = 36'hf5dee748f;
            11'd184: table_out = 36'hf5e123f5d;
            11'd185: table_out = 36'hf5e3606b4;
            11'd186: table_out = 36'hf5e59ca93;
            11'd187: table_out = 36'hf5e7d8afc;
            11'd188: table_out = 36'hf5ea147ef;
            11'd189: table_out = 36'hf5ec5016e;
            11'd190: table_out = 36'hf5ee8b778;
            11'd191: table_out = 36'hf5f0c6a0f;
            11'd192: table_out = 36'hf5f301932;
            11'd193: table_out = 36'hf5f53c4e3;
            11'd194: table_out = 36'hf5f776d23;
            11'd195: table_out = 36'hf5f9b11f2;
            11'd196: table_out = 36'hf5fbeb350;
            11'd197: table_out = 36'hf5fe2513f;
            11'd198: table_out = 36'hf6005ebbf;
            11'd199: table_out = 36'hf602982d0;
            11'd200: table_out = 36'hf604d1674;
            11'd201: table_out = 36'hf6070a6ab;
            11'd202: table_out = 36'hf60943375;
            11'd203: table_out = 36'hf60b7bcd4;
            11'd204: table_out = 36'hf60db42c8;
            11'd205: table_out = 36'hf60fec551;
            11'd206: table_out = 36'hf61224471;
            11'd207: table_out = 36'hf6145c028;
            11'd208: table_out = 36'hf61693876;
            11'd209: table_out = 36'hf618cad5d;
            11'd210: table_out = 36'hf61b01edc;
            11'd211: table_out = 36'hf61d38cf5;
            11'd212: table_out = 36'hf61f6f7a9;
            11'd213: table_out = 36'hf621a5ef7;
            11'd214: table_out = 36'hf623dc2e1;
            11'd215: table_out = 36'hf62612366;
            11'd216: table_out = 36'hf62848089;
            11'd217: table_out = 36'hf62a7da49;
            11'd218: table_out = 36'hf62cb30a8;
            11'd219: table_out = 36'hf62ee83a5;
            11'd220: table_out = 36'hf6311d341;
            11'd221: table_out = 36'hf63351f7e;
            11'd222: table_out = 36'hf6358685b;
            11'd223: table_out = 36'hf637badda;
            11'd224: table_out = 36'hf639eeffa;
            11'd225: table_out = 36'hf63c22ebe;
            11'd226: table_out = 36'hf63e56a24;
            11'd227: table_out = 36'hf6408a22f;
            11'd228: table_out = 36'hf642bd6de;
            11'd229: table_out = 36'hf644f0832;
            11'd230: table_out = 36'hf6472362c;
            11'd231: table_out = 36'hf649560cc;
            11'd232: table_out = 36'hf64b88814;
            11'd233: table_out = 36'hf64dbac03;
            11'd234: table_out = 36'hf64fecc9b;
            11'd235: table_out = 36'hf6521e9dc;
            11'd236: table_out = 36'hf654503c7;
            11'd237: table_out = 36'hf65681a5b;
            11'd238: table_out = 36'hf658b2d9b;
            11'd239: table_out = 36'hf65ae3d86;
            11'd240: table_out = 36'hf65d14a1e;
            11'd241: table_out = 36'hf65f45362;
            11'd242: table_out = 36'hf66175954;
            11'd243: table_out = 36'hf663a5bf3;
            11'd244: table_out = 36'hf665d5b42;
            11'd245: table_out = 36'hf66805740;
            11'd246: table_out = 36'hf66a34fee;
            11'd247: table_out = 36'hf66c6454c;
            11'd248: table_out = 36'hf66e9375c;
            11'd249: table_out = 36'hf670c261d;
            11'd250: table_out = 36'hf672f1191;
            11'd251: table_out = 36'hf6751f9b8;
            11'd252: table_out = 36'hf6774de93;
            11'd253: table_out = 36'hf6797c022;
            11'd254: table_out = 36'hf67ba9e66;
            11'd255: table_out = 36'hf67dd7960;
            11'd256: table_out = 36'hf68005110;
            11'd257: table_out = 36'hf68232576;
            11'd258: table_out = 36'hf6845f694;
            11'd259: table_out = 36'hf6868c46b;
            11'd260: table_out = 36'hf688b8efa;
            11'd261: table_out = 36'hf68ae5642;
            11'd262: table_out = 36'hf68d11a44;
            11'd263: table_out = 36'hf68f3db00;
            11'd264: table_out = 36'hf69169878;
            11'd265: table_out = 36'hf693952ac;
            11'd266: table_out = 36'hf695c099c;
            11'd267: table_out = 36'hf697ebd49;
            11'd268: table_out = 36'hf69a16db3;
            11'd269: table_out = 36'hf69c41adc;
            11'd270: table_out = 36'hf69e6c4c4;
            11'd271: table_out = 36'hf6a096b6b;
            11'd272: table_out = 36'hf6a2c0ed2;
            11'd273: table_out = 36'hf6a4eaef9;
            11'd274: table_out = 36'hf6a714be3;
            11'd275: table_out = 36'hf6a93e58d;
            11'd276: table_out = 36'hf6ab67bfb;
            11'd277: table_out = 36'hf6ad90f2b;
            11'd278: table_out = 36'hf6afb9f1f;
            11'd279: table_out = 36'hf6b1e2bd8;
            11'd280: table_out = 36'hf6b40b555;
            11'd281: table_out = 36'hf6b633b98;
            11'd282: table_out = 36'hf6b85bea1;
            11'd283: table_out = 36'hf6ba83e71;
            11'd284: table_out = 36'hf6bcabb08;
            11'd285: table_out = 36'hf6bed3467;
            11'd286: table_out = 36'hf6c0faa8e;
            11'd287: table_out = 36'hf6c321d7f;
            11'd288: table_out = 36'hf6c548d39;
            11'd289: table_out = 36'hf6c76f9be;
            11'd290: table_out = 36'hf6c99630d;
            11'd291: table_out = 36'hf6cbbc928;
            11'd292: table_out = 36'hf6cde2c0f;
            11'd293: table_out = 36'hf6d008bc3;
            11'd294: table_out = 36'hf6d22e844;
            11'd295: table_out = 36'hf6d454193;
            11'd296: table_out = 36'hf6d6797b1;
            11'd297: table_out = 36'hf6d89ea9e;
            11'd298: table_out = 36'hf6dac3a5a;
            11'd299: table_out = 36'hf6dce86e6;
            11'd300: table_out = 36'hf6df0d044;
            11'd301: table_out = 36'hf6e131673;
            11'd302: table_out = 36'hf6e355974;
            11'd303: table_out = 36'hf6e579947;
            11'd304: table_out = 36'hf6e79d5ee;
            11'd305: table_out = 36'hf6e9c0f69;
            11'd306: table_out = 36'hf6ebe45b8;
            11'd307: table_out = 36'hf6ee078dc;
            11'd308: table_out = 36'hf6f02a8d5;
            11'd309: table_out = 36'hf6f24d5a5;
            11'd310: table_out = 36'hf6f46ff4b;
            11'd311: table_out = 36'hf6f6925c9;
            11'd312: table_out = 36'hf6f8b491f;
            11'd313: table_out = 36'hf6fad694d;
            11'd314: table_out = 36'hf6fcf8654;
            11'd315: table_out = 36'hf6ff1a035;
            11'd316: table_out = 36'hf7013b6f0;
            11'd317: table_out = 36'hf7035ca86;
            11'd318: table_out = 36'hf7057daf8;
            11'd319: table_out = 36'hf7079e845;
            11'd320: table_out = 36'hf709bf26f;
            11'd321: table_out = 36'hf70bdf976;
            11'd322: table_out = 36'hf70dffd5b;
            11'd323: table_out = 36'hf7101fe1e;
            11'd324: table_out = 36'hf7123fbc0;
            11'd325: table_out = 36'hf7145f641;
            11'd326: table_out = 36'hf7167eda3;
            11'd327: table_out = 36'hf7189e1e5;
            11'd328: table_out = 36'hf71abd308;
            11'd329: table_out = 36'hf71cdc10d;
            11'd330: table_out = 36'hf71efabf4;
            11'd331: table_out = 36'hf721193be;
            11'd332: table_out = 36'hf7233786c;
            11'd333: table_out = 36'hf725559fd;
            11'd334: table_out = 36'hf72773873;
            11'd335: table_out = 36'hf729913cf;
            11'd336: table_out = 36'hf72baec10;
            11'd337: table_out = 36'hf72dcc137;
            11'd338: table_out = 36'hf72fe9346;
            11'd339: table_out = 36'hf7320623b;
            11'd340: table_out = 36'hf73422e19;
            11'd341: table_out = 36'hf7363f6e0;
            11'd342: table_out = 36'hf7385bc8f;
            11'd343: table_out = 36'hf73a77f28;
            11'd344: table_out = 36'hf73c93eac;
            11'd345: table_out = 36'hf73eafb1a;
            11'd346: table_out = 36'hf740cb474;
            11'd347: table_out = 36'hf742e6ab9;
            11'd348: table_out = 36'hf74501deb;
            11'd349: table_out = 36'hf7471ce0b;
            11'd350: table_out = 36'hf74937b17;
            11'd351: table_out = 36'hf74b52512;
            11'd352: table_out = 36'hf74d6cbfc;
            11'd353: table_out = 36'hf74f86fd5;
            11'd354: table_out = 36'hf751a109e;
            11'd355: table_out = 36'hf753bae58;
            11'd356: table_out = 36'hf755d4902;
            11'd357: table_out = 36'hf757ee09e;
            11'd358: table_out = 36'hf75a0752c;
            11'd359: table_out = 36'hf75c206ad;
            11'd360: table_out = 36'hf75e39521;
            11'd361: table_out = 36'hf76052089;
            11'd362: table_out = 36'hf7626a8e5;
            11'd363: table_out = 36'hf76482e36;
            11'd364: table_out = 36'hf7669b07c;
            11'd365: table_out = 36'hf768b2fb9;
            11'd366: table_out = 36'hf76acabec;
            11'd367: table_out = 36'hf76ce2516;
            11'd368: table_out = 36'hf76ef9b37;
            11'd369: table_out = 36'hf77110e51;
            11'd370: table_out = 36'hf77327e63;
            11'd371: table_out = 36'hf7753eb6f;
            11'd372: table_out = 36'hf77755575;
            11'd373: table_out = 36'hf7796bc75;
            11'd374: table_out = 36'hf77b82070;
            11'd375: table_out = 36'hf77d98166;
            11'd376: table_out = 36'hf77fadf58;
            11'd377: table_out = 36'hf781c3a47;
            11'd378: table_out = 36'hf783d9233;
            11'd379: table_out = 36'hf785ee71d;
            11'd380: table_out = 36'hf78803905;
            11'd381: table_out = 36'hf78a187eb;
            11'd382: table_out = 36'hf78c2d3d1;
            11'd383: table_out = 36'hf78e41cb7;
            11'd384: table_out = 36'hf7905629d;
            11'd385: table_out = 36'hf7926a584;
            11'd386: table_out = 36'hf7947e56c;
            11'd387: table_out = 36'hf79692256;
            11'd388: table_out = 36'hf798a5c43;
            11'd389: table_out = 36'hf79ab9333;
            11'd390: table_out = 36'hf79ccc726;
            11'd391: table_out = 36'hf79edf81e;
            11'd392: table_out = 36'hf7a0f261a;
            11'd393: table_out = 36'hf7a30511b;
            11'd394: table_out = 36'hf7a517922;
            11'd395: table_out = 36'hf7a729e30;
            11'd396: table_out = 36'hf7a93c044;
            11'd397: table_out = 36'hf7ab4df5f;
            11'd398: table_out = 36'hf7ad5fb83;
            11'd399: table_out = 36'hf7af714af;
            11'd400: table_out = 36'hf7b182ae3;
            11'd401: table_out = 36'hf7b393e21;
            11'd402: table_out = 36'hf7b5a4e69;
            11'd403: table_out = 36'hf7b7b5bbc;
            11'd404: table_out = 36'hf7b9c661a;
            11'd405: table_out = 36'hf7bbd6d83;
            11'd406: table_out = 36'hf7bde71f8;
            11'd407: table_out = 36'hf7bff737a;
            11'd408: table_out = 36'hf7c207209;
            11'd409: table_out = 36'hf7c416da6;
            11'd410: table_out = 36'hf7c626651;
            11'd411: table_out = 36'hf7c835c0b;
            11'd412: table_out = 36'hf7ca44ed4;
            11'd413: table_out = 36'hf7cc53ead;
            11'd414: table_out = 36'hf7ce62b96;
            11'd415: table_out = 36'hf7d071590;
            11'd416: table_out = 36'hf7d27fc9b;
            11'd417: table_out = 36'hf7d48e0b8;
            11'd418: table_out = 36'hf7d69c1e8;
            11'd419: table_out = 36'hf7d8aa02a;
            11'd420: table_out = 36'hf7dab7b80;
            11'd421: table_out = 36'hf7dcc53ea;
            11'd422: table_out = 36'hf7ded2968;
            11'd423: table_out = 36'hf7e0dfbfc;
            11'd424: table_out = 36'hf7e2ecba5;
            11'd425: table_out = 36'hf7e4f9863;
            11'd426: table_out = 36'hf7e706239;
            11'd427: table_out = 36'hf7e912925;
            11'd428: table_out = 36'hf7eb1ed2a;
            11'd429: table_out = 36'hf7ed2ae46;
            11'd430: table_out = 36'hf7ef36c7b;
            11'd431: table_out = 36'hf7f1427c9;
            11'd432: table_out = 36'hf7f34e030;
            11'd433: table_out = 36'hf7f5595b2;
            11'd434: table_out = 36'hf7f76484e;
            11'd435: table_out = 36'hf7f96f806;
            11'd436: table_out = 36'hf7fb7a4d9;
            11'd437: table_out = 36'hf7fd84ec9;
            11'd438: table_out = 36'hf7ff8f5d5;
            11'd439: table_out = 36'hf801999ff;
            11'd440: table_out = 36'hf803a3b46;
            11'd441: table_out = 36'hf805ad9ab;
            11'd442: table_out = 36'hf807b7530;
            11'd443: table_out = 36'hf809c0dd3;
            11'd444: table_out = 36'hf80bca396;
            11'd445: table_out = 36'hf80dd367a;
            11'd446: table_out = 36'hf80fdc67e;
            11'd447: table_out = 36'hf811e53a4;
            11'd448: table_out = 36'hf813eddeb;
            11'd449: table_out = 36'hf815f6555;
            11'd450: table_out = 36'hf817fe9e2;
            11'd451: table_out = 36'hf81a06b92;
            11'd452: table_out = 36'hf81c0ea65;
            11'd453: table_out = 36'hf81e1665d;
            11'd454: table_out = 36'hf8201df7a;
            11'd455: table_out = 36'hf822255bc;
            11'd456: table_out = 36'hf8242c924;
            11'd457: table_out = 36'hf826339b3;
            11'd458: table_out = 36'hf8283a768;
            11'd459: table_out = 36'hf82a41244;
            11'd460: table_out = 36'hf82c47a48;
            11'd461: table_out = 36'hf82e4df75;
            11'd462: table_out = 36'hf830541cb;
            11'd463: table_out = 36'hf8325a149;
            11'd464: table_out = 36'hf8345fdf2;
            11'd465: table_out = 36'hf836657c5;
            11'd466: table_out = 36'hf8386aec3;
            11'd467: table_out = 36'hf83a702ec;
            11'd468: table_out = 36'hf83c75440;
            11'd469: table_out = 36'hf83e7a2c2;
            11'd470: table_out = 36'hf8407ee70;
            11'd471: table_out = 36'hf8428374b;
            11'd472: table_out = 36'hf84487d54;
            11'd473: table_out = 36'hf8468c08b;
            11'd474: table_out = 36'hf848900f1;
            11'd475: table_out = 36'hf84a93e87;
            11'd476: table_out = 36'hf84c9794c;
            11'd477: table_out = 36'hf84e9b141;
            11'd478: table_out = 36'hf8509e667;
            11'd479: table_out = 36'hf852a18be;
            11'd480: table_out = 36'hf854a4847;
            11'd481: table_out = 36'hf856a7502;
            11'd482: table_out = 36'hf858a9ef0;
            11'd483: table_out = 36'hf85aac611;
            11'd484: table_out = 36'hf85caea66;
            11'd485: table_out = 36'hf85eb0bef;
            11'd486: table_out = 36'hf860b2aac;
            11'd487: table_out = 36'hf862b469f;
            11'd488: table_out = 36'hf864b5fc7;
            11'd489: table_out = 36'hf866b7626;
            11'd490: table_out = 36'hf868b89bb;
            11'd491: table_out = 36'hf86ab9a86;
            11'd492: table_out = 36'hf86cba88a;
            11'd493: table_out = 36'hf86ebb3c6;
            11'd494: table_out = 36'hf870bbc3a;
            11'd495: table_out = 36'hf872bc1e7;
            11'd496: table_out = 36'hf874bc4cd;
            11'd497: table_out = 36'hf876bc4ee;
            11'd498: table_out = 36'hf878bc249;
            11'd499: table_out = 36'hf87abbcde;
            11'd500: table_out = 36'hf87cbb4b0;
            11'd501: table_out = 36'hf87eba9bd;
            11'd502: table_out = 36'hf880b9c06;
            11'd503: table_out = 36'hf882b8b8c;
            11'd504: table_out = 36'hf884b7850;
            11'd505: table_out = 36'hf886b6251;
            11'd506: table_out = 36'hf888b4991;
            11'd507: table_out = 36'hf88ab2e0f;
            11'd508: table_out = 36'hf88cb0fcd;
            11'd509: table_out = 36'hf88eaeeca;
            11'd510: table_out = 36'hf890acb08;
            11'd511: table_out = 36'hf892aa486;
            11'd512: table_out = 36'hf894a7b45;
            11'd513: table_out = 36'hf896a4f46;
            11'd514: table_out = 36'hf898a2088;
            11'd515: table_out = 36'hf89a9ef0e;
            11'd516: table_out = 36'hf89c9bad6;
            11'd517: table_out = 36'hf89e983e2;
            11'd518: table_out = 36'hf8a094a32;
            11'd519: table_out = 36'hf8a290dc6;
            11'd520: table_out = 36'hf8a48ce9f;
            11'd521: table_out = 36'hf8a688cbd;
            11'd522: table_out = 36'hf8a884822;
            11'd523: table_out = 36'hf8aa800cc;
            11'd524: table_out = 36'hf8ac7b6be;
            11'd525: table_out = 36'hf8ae769f6;
            11'd526: table_out = 36'hf8b071a76;
            11'd527: table_out = 36'hf8b26c83f;
            11'd528: table_out = 36'hf8b467350;
            11'd529: table_out = 36'hf8b661baa;
            11'd530: table_out = 36'hf8b85c14d;
            11'd531: table_out = 36'hf8ba5643b;
            11'd532: table_out = 36'hf8bc50473;
            11'd533: table_out = 36'hf8be4a1f6;
            11'd534: table_out = 36'hf8c043cc5;
            11'd535: table_out = 36'hf8c23d4df;
            11'd536: table_out = 36'hf8c436a46;
            11'd537: table_out = 36'hf8c62fcf9;
            11'd538: table_out = 36'hf8c828cfa;
            11'd539: table_out = 36'hf8ca21a49;
            11'd540: table_out = 36'hf8cc1a4e5;
            11'd541: table_out = 36'hf8ce12cd1;
            11'd542: table_out = 36'hf8d00b20b;
            11'd543: table_out = 36'hf8d203495;
            11'd544: table_out = 36'hf8d3fb46f;
            11'd545: table_out = 36'hf8d5f319a;
            11'd546: table_out = 36'hf8d7eac15;
            11'd547: table_out = 36'hf8d9e23e2;
            11'd548: table_out = 36'hf8dbd9901;
            11'd549: table_out = 36'hf8ddd0b72;
            11'd550: table_out = 36'hf8dfc7b36;
            11'd551: table_out = 36'hf8e1be84c;
            11'd552: table_out = 36'hf8e3b52b7;
            11'd553: table_out = 36'hf8e5aba76;
            11'd554: table_out = 36'hf8e7a1f89;
            11'd555: table_out = 36'hf8e9981f2;
            11'd556: table_out = 36'hf8eb8e1b0;
            11'd557: table_out = 36'hf8ed83ec3;
            11'd558: table_out = 36'hf8ef7992e;
            11'd559: table_out = 36'hf8f16f0ef;
            11'd560: table_out = 36'hf8f364607;
            11'd561: table_out = 36'hf8f559877;
            11'd562: table_out = 36'hf8f74e840;
            11'd563: table_out = 36'hf8f943561;
            11'd564: table_out = 36'hf8fb37fdb;
            11'd565: table_out = 36'hf8fd2c7ae;
            11'd566: table_out = 36'hf8ff20cdc;
            11'd567: table_out = 36'hf90114f64;
            11'd568: table_out = 36'hf90308f47;
            11'd569: table_out = 36'hf904fcc85;
            11'd570: table_out = 36'hf906f071f;
            11'd571: table_out = 36'hf908e3f16;
            11'd572: table_out = 36'hf90ad7469;
            11'd573: table_out = 36'hf90cca719;
            11'd574: table_out = 36'hf90ebd726;
            11'd575: table_out = 36'hf910b0492;
            11'd576: table_out = 36'hf912a2f5c;
            11'd577: table_out = 36'hf91495785;
            11'd578: table_out = 36'hf91687d0e;
            11'd579: table_out = 36'hf91879ff6;
            11'd580: table_out = 36'hf91a6c03e;
            11'd581: table_out = 36'hf91c5dde8;
            11'd582: table_out = 36'hf91e4f8f2;
            11'd583: table_out = 36'hf9204115e;
            11'd584: table_out = 36'hf9223272b;
            11'd585: table_out = 36'hf92423a5c;
            11'd586: table_out = 36'hf92614aef;
            11'd587: table_out = 36'hf928058e5;
            11'd588: table_out = 36'hf929f6440;
            11'd589: table_out = 36'hf92be6cfe;
            11'd590: table_out = 36'hf92dd7321;
            11'd591: table_out = 36'hf92fc76a9;
            11'd592: table_out = 36'hf931b7797;
            11'd593: table_out = 36'hf933a75ea;
            11'd594: table_out = 36'hf935971a4;
            11'd595: table_out = 36'hf93786ac5;
            11'd596: table_out = 36'hf9397614d;
            11'd597: table_out = 36'hf93b6553d;
            11'd598: table_out = 36'hf93d54695;
            11'd599: table_out = 36'hf93f43555;
            11'd600: table_out = 36'hf9413217f;
            11'd601: table_out = 36'hf94320b11;
            11'd602: table_out = 36'hf9450f20e;
            11'd603: table_out = 36'hf946fd675;
            11'd604: table_out = 36'hf948eb847;
            11'd605: table_out = 36'hf94ad9784;
            11'd606: table_out = 36'hf94cc742c;
            11'd607: table_out = 36'hf94eb4e41;
            11'd608: table_out = 36'hf950a25c2;
            11'd609: table_out = 36'hf9528faaf;
            11'd610: table_out = 36'hf9547cd0b;
            11'd611: table_out = 36'hf95669cd3;
            11'd612: table_out = 36'hf95856a0a;
            11'd613: table_out = 36'hf95a434b0;
            11'd614: table_out = 36'hf95c2fcc5;
            11'd615: table_out = 36'hf95e1c249;
            11'd616: table_out = 36'hf9600853d;
            11'd617: table_out = 36'hf961f45a1;
            11'd618: table_out = 36'hf963e0376;
            11'd619: table_out = 36'hf965cbebc;
            11'd620: table_out = 36'hf967b7774;
            11'd621: table_out = 36'hf969a2d9e;
            11'd622: table_out = 36'hf96b8e13a;
            11'd623: table_out = 36'hf96d79249;
            11'd624: table_out = 36'hf96f640cc;
            11'd625: table_out = 36'hf9714ecc2;
            11'd626: table_out = 36'hf9733962c;
            11'd627: table_out = 36'hf97523d0b;
            11'd628: table_out = 36'hf9770e15f;
            11'd629: table_out = 36'hf978f8328;
            11'd630: table_out = 36'hf97ae2267;
            11'd631: table_out = 36'hf97ccbf1c;
            11'd632: table_out = 36'hf97eb5948;
            11'd633: table_out = 36'hf9809f0eb;
            11'd634: table_out = 36'hf98288605;
            11'd635: table_out = 36'hf98471897;
            11'd636: table_out = 36'hf9865a8a2;
            11'd637: table_out = 36'hf98843626;
            11'd638: table_out = 36'hf98a2c122;
            11'd639: table_out = 36'hf98c14998;
            11'd640: table_out = 36'hf98dfcf89;
            11'd641: table_out = 36'hf98fe52f3;
            11'd642: table_out = 36'hf991cd3d9;
            11'd643: table_out = 36'hf993b523a;
            11'd644: table_out = 36'hf9959ce16;
            11'd645: table_out = 36'hf9978476f;
            11'd646: table_out = 36'hf9996be44;
            11'd647: table_out = 36'hf99b53296;
            11'd648: table_out = 36'hf99d3a465;
            11'd649: table_out = 36'hf99f213b2;
            11'd650: table_out = 36'hf9a10807d;
            11'd651: table_out = 36'hf9a2eeac7;
            11'd652: table_out = 36'hf9a4d5290;
            11'd653: table_out = 36'hf9a6bb7d8;
            11'd654: table_out = 36'hf9a8a1aa0;
            11'd655: table_out = 36'hf9aa87ae8;
            11'd656: table_out = 36'hf9ac6d8b1;
            11'd657: table_out = 36'hf9ae533fb;
            11'd658: table_out = 36'hf9b038cc6;
            11'd659: table_out = 36'hf9b21e313;
            11'd660: table_out = 36'hf9b4036e3;
            11'd661: table_out = 36'hf9b5e8835;
            11'd662: table_out = 36'hf9b7cd70a;
            11'd663: table_out = 36'hf9b9b2363;
            11'd664: table_out = 36'hf9bb96d3f;
            11'd665: table_out = 36'hf9bd7b4a0;
            11'd666: table_out = 36'hf9bf5f986;
            11'd667: table_out = 36'hf9c143bf1;
            11'd668: table_out = 36'hf9c327be1;
            11'd669: table_out = 36'hf9c50b957;
            11'd670: table_out = 36'hf9c6ef454;
            11'd671: table_out = 36'hf9c8d2cd7;
            11'd672: table_out = 36'hf9cab62e2;
            11'd673: table_out = 36'hf9cc99674;
            11'd674: table_out = 36'hf9ce7c78e;
            11'd675: table_out = 36'hf9d05f630;
            11'd676: table_out = 36'hf9d24225c;
            11'd677: table_out = 36'hf9d424c10;
            11'd678: table_out = 36'hf9d60734e;
            11'd679: table_out = 36'hf9d7e9816;
            11'd680: table_out = 36'hf9d9cba68;
            11'd681: table_out = 36'hf9dbada45;
            11'd682: table_out = 36'hf9dd8f7ad;
            11'd683: table_out = 36'hf9df712a1;
            11'd684: table_out = 36'hf9e152b21;
            11'd685: table_out = 36'hf9e33412d;
            11'd686: table_out = 36'hf9e5154c6;
            11'd687: table_out = 36'hf9e6f65ec;
            11'd688: table_out = 36'hf9e8d74a0;
            11'd689: table_out = 36'hf9eab80e2;
            11'd690: table_out = 36'hf9ec98ab2;
            11'd691: table_out = 36'hf9ee79211;
            11'd692: table_out = 36'hf9f0596ff;
            11'd693: table_out = 36'hf9f23997c;
            11'd694: table_out = 36'hf9f41998a;
            11'd695: table_out = 36'hf9f5f9728;
            11'd696: table_out = 36'hf9f7d9256;
            11'd697: table_out = 36'hf9f9b8b16;
            11'd698: table_out = 36'hf9fb98168;
            11'd699: table_out = 36'hf9fd7754b;
            11'd700: table_out = 36'hf9ff566c0;
            11'd701: table_out = 36'hfa01355c9;
            11'd702: table_out = 36'hfa0314264;
            11'd703: table_out = 36'hfa04f2c93;
            11'd704: table_out = 36'hfa06d1456;
            11'd705: table_out = 36'hfa08af9ad;
            11'd706: table_out = 36'hfa0a8dc99;
            11'd707: table_out = 36'hfa0c6bd1a;
            11'd708: table_out = 36'hfa0e49b30;
            11'd709: table_out = 36'hfa10276dd;
            11'd710: table_out = 36'hfa120501f;
            11'd711: table_out = 36'hfa13e26f8;
            11'd712: table_out = 36'hfa15bfb68;
            11'd713: table_out = 36'hfa179cd70;
            11'd714: table_out = 36'hfa1979d0f;
            11'd715: table_out = 36'hfa1b56a47;
            11'd716: table_out = 36'hfa1d33517;
            11'd717: table_out = 36'hfa1f0fd80;
            11'd718: table_out = 36'hfa20ec383;
            11'd719: table_out = 36'hfa22c871f;
            11'd720: table_out = 36'hfa24a4856;
            11'd721: table_out = 36'hfa2680726;
            11'd722: table_out = 36'hfa285c392;
            11'd723: table_out = 36'hfa2a37d99;
            11'd724: table_out = 36'hfa2c1353c;
            11'd725: table_out = 36'hfa2deea7b;
            11'd726: table_out = 36'hfa2fc9d56;
            11'd727: table_out = 36'hfa31a4dce;
            11'd728: table_out = 36'hfa337fbe4;
            11'd729: table_out = 36'hfa355a797;
            11'd730: table_out = 36'hfa37350e8;
            11'd731: table_out = 36'hfa390f7d7;
            11'd732: table_out = 36'hfa3ae9c65;
            11'd733: table_out = 36'hfa3cc3e92;
            11'd734: table_out = 36'hfa3e9de5f;
            11'd735: table_out = 36'hfa4077bcb;
            11'd736: table_out = 36'hfa42516d8;
            11'd737: table_out = 36'hfa442af85;
            11'd738: table_out = 36'hfa46045d4;
            11'd739: table_out = 36'hfa47dd9c4;
            11'd740: table_out = 36'hfa49b6b55;
            11'd741: table_out = 36'hfa4b8fa89;
            11'd742: table_out = 36'hfa4d68760;
            11'd743: table_out = 36'hfa4f411d9;
            11'd744: table_out = 36'hfa51199f6;
            11'd745: table_out = 36'hfa52f1fb6;
            11'd746: table_out = 36'hfa54ca31a;
            11'd747: table_out = 36'hfa56a2423;
            11'd748: table_out = 36'hfa587a2d1;
            11'd749: table_out = 36'hfa5a51f23;
            11'd750: table_out = 36'hfa5c2991c;
            11'd751: table_out = 36'hfa5e010ba;
            11'd752: table_out = 36'hfa5fd85ff;
            11'd753: table_out = 36'hfa61af8ea;
            11'd754: table_out = 36'hfa638697c;
            11'd755: table_out = 36'hfa655d7b6;
            11'd756: table_out = 36'hfa6734398;
            11'd757: table_out = 36'hfa690ad22;
            11'd758: table_out = 36'hfa6ae1454;
            11'd759: table_out = 36'hfa6cb792f;
            11'd760: table_out = 36'hfa6e8dbb4;
            11'd761: table_out = 36'hfa7063be2;
            11'd762: table_out = 36'hfa72399ba;
            11'd763: table_out = 36'hfa740f53d;
            11'd764: table_out = 36'hfa75e4e6b;
            11'd765: table_out = 36'hfa77ba543;
            11'd766: table_out = 36'hfa798f9c8;
            11'd767: table_out = 36'hfa7b64bf8;
            11'd768: table_out = 36'hfa7d39bd4;
            11'd769: table_out = 36'hfa7f0e95d;
            11'd770: table_out = 36'hfa80e3493;
            11'd771: table_out = 36'hfa82b7d77;
            11'd772: table_out = 36'hfa848c408;
            11'd773: table_out = 36'hfa8660847;
            11'd774: table_out = 36'hfa8834a35;
            11'd775: table_out = 36'hfa8a089d1;
            11'd776: table_out = 36'hfa8bdc71d;
            11'd777: table_out = 36'hfa8db0219;
            11'd778: table_out = 36'hfa8f83ac4;
            11'd779: table_out = 36'hfa915711f;
            11'd780: table_out = 36'hfa932a52c;
            11'd781: table_out = 36'hfa94fd6e9;
            11'd782: table_out = 36'hfa96d0658;
            11'd783: table_out = 36'hfa98a3378;
            11'd784: table_out = 36'hfa9a75e4b;
            11'd785: table_out = 36'hfa9c486d0;
            11'd786: table_out = 36'hfa9e1ad08;
            11'd787: table_out = 36'hfa9fed0f4;
            11'd788: table_out = 36'hfaa1bf293;
            11'd789: table_out = 36'hfaa3911e5;
            11'd790: table_out = 36'hfaa562eed;
            11'd791: table_out = 36'hfaa7349a8;
            11'd792: table_out = 36'hfaa906219;
            11'd793: table_out = 36'hfaaad783f;
            11'd794: table_out = 36'hfaaca8c1b;
            11'd795: table_out = 36'hfaae79dae;
            11'd796: table_out = 36'hfab04acf6;
            11'd797: table_out = 36'hfab21b9f6;
            11'd798: table_out = 36'hfab3ec4ac;
            11'd799: table_out = 36'hfab5bcd1a;
            11'd800: table_out = 36'hfab78d341;
            11'd801: table_out = 36'hfab95d71f;
            11'd802: table_out = 36'hfabb2d8b6;
            11'd803: table_out = 36'hfabcfd806;
            11'd804: table_out = 36'hfabecd50f;
            11'd805: table_out = 36'hfac09cfd3;
            11'd806: table_out = 36'hfac26c850;
            11'd807: table_out = 36'hfac43be87;
            11'd808: table_out = 36'hfac60b27a;
            11'd809: table_out = 36'hfac7da427;
            11'd810: table_out = 36'hfac9a9390;
            11'd811: table_out = 36'hfacb780b5;
            11'd812: table_out = 36'hfacd46b96;
            11'd813: table_out = 36'hfacf15433;
            11'd814: table_out = 36'hfad0e3a8e;
            11'd815: table_out = 36'hfad2b1ea6;
            11'd816: table_out = 36'hfad48007b;
            11'd817: table_out = 36'hfad64e00e;
            11'd818: table_out = 36'hfad81bd60;
            11'd819: table_out = 36'hfad9e9870;
            11'd820: table_out = 36'hfadbb713f;
            11'd821: table_out = 36'hfadd847ce;
            11'd822: table_out = 36'hfadf51c1d;
            11'd823: table_out = 36'hfae11ee2b;
            11'd824: table_out = 36'hfae2ebdfa;
            11'd825: table_out = 36'hfae4b8b8a;
            11'd826: table_out = 36'hfae6856db;
            11'd827: table_out = 36'hfae851fed;
            11'd828: table_out = 36'hfaea1e6c1;
            11'd829: table_out = 36'hfaebeab58;
            11'd830: table_out = 36'hfaedb6db0;
            11'd831: table_out = 36'hfaef82dcc;
            11'd832: table_out = 36'hfaf14ebab;
            11'd833: table_out = 36'hfaf31a74e;
            11'd834: table_out = 36'hfaf4e60b4;
            11'd835: table_out = 36'hfaf6b17df;
            11'd836: table_out = 36'hfaf87ccce;
            11'd837: table_out = 36'hfafa47f83;
            11'd838: table_out = 36'hfafc12ffc;
            11'd839: table_out = 36'hfafddde3c;
            11'd840: table_out = 36'hfaffa8a41;
            11'd841: table_out = 36'hfb017340d;
            11'd842: table_out = 36'hfb033db9f;
            11'd843: table_out = 36'hfb05080f9;
            11'd844: table_out = 36'hfb06d2419;
            11'd845: table_out = 36'hfb089c502;
            11'd846: table_out = 36'hfb0a663b2;
            11'd847: table_out = 36'hfb0c3002b;
            11'd848: table_out = 36'hfb0df9a6d;
            11'd849: table_out = 36'hfb0fc3278;
            11'd850: table_out = 36'hfb118c84c;
            11'd851: table_out = 36'hfb1355beb;
            11'd852: table_out = 36'hfb151ed53;
            11'd853: table_out = 36'hfb16e7c85;
            11'd854: table_out = 36'hfb18b0983;
            11'd855: table_out = 36'hfb1a7944c;
            11'd856: table_out = 36'hfb1c41ce0;
            11'd857: table_out = 36'hfb1e0a340;
            11'd858: table_out = 36'hfb1fd276c;
            11'd859: table_out = 36'hfb219a965;
            11'd860: table_out = 36'hfb236292a;
            11'd861: table_out = 36'hfb252a6bd;
            11'd862: table_out = 36'hfb26f221d;
            11'd863: table_out = 36'hfb28b9b4c;
            11'd864: table_out = 36'hfb2a81248;
            11'd865: table_out = 36'hfb2c48713;
            11'd866: table_out = 36'hfb2e0f9ad;
            11'd867: table_out = 36'hfb2fd6a16;
            11'd868: table_out = 36'hfb319d84e;
            11'd869: table_out = 36'hfb3364457;
            11'd870: table_out = 36'hfb352ae30;
            11'd871: table_out = 36'hfb36f15d9;
            11'd872: table_out = 36'hfb38b7b53;
            11'd873: table_out = 36'hfb3a7de9f;
            11'd874: table_out = 36'hfb3c43fbc;
            11'd875: table_out = 36'hfb3e09eab;
            11'd876: table_out = 36'hfb3fcfb6c;
            11'd877: table_out = 36'hfb4195600;
            11'd878: table_out = 36'hfb435ae66;
            11'd879: table_out = 36'hfb45204a0;
            11'd880: table_out = 36'hfb46e58ae;
            11'd881: table_out = 36'hfb48aaa8f;
            11'd882: table_out = 36'hfb4a6fa45;
            11'd883: table_out = 36'hfb4c347cf;
            11'd884: table_out = 36'hfb4df932f;
            11'd885: table_out = 36'hfb4fbdc63;
            11'd886: table_out = 36'hfb518236d;
            11'd887: table_out = 36'hfb534684d;
            11'd888: table_out = 36'hfb550ab03;
            11'd889: table_out = 36'hfb56ceb90;
            11'd890: table_out = 36'hfb58929f4;
            11'd891: table_out = 36'hfb5a5662f;
            11'd892: table_out = 36'hfb5c1a041;
            11'd893: table_out = 36'hfb5ddd82c;
            11'd894: table_out = 36'hfb5fa0dee;
            11'd895: table_out = 36'hfb616418a;
            11'd896: table_out = 36'hfb63272fe;
            11'd897: table_out = 36'hfb64ea24b;
            11'd898: table_out = 36'hfb66acf72;
            11'd899: table_out = 36'hfb686fa73;
            11'd900: table_out = 36'hfb6a3234d;
            11'd901: table_out = 36'hfb6bf4a03;
            11'd902: table_out = 36'hfb6db6e93;
            11'd903: table_out = 36'hfb6f790ff;
            11'd904: table_out = 36'hfb713b146;
            11'd905: table_out = 36'hfb72fcf68;
            11'd906: table_out = 36'hfb74beb67;
            11'd907: table_out = 36'hfb7680543;
            11'd908: table_out = 36'hfb7841cfb;
            11'd909: table_out = 36'hfb7a03290;
            11'd910: table_out = 36'hfb7bc4603;
            11'd911: table_out = 36'hfb7d85754;
            11'd912: table_out = 36'hfb7f46682;
            11'd913: table_out = 36'hfb8107390;
            11'd914: table_out = 36'hfb82c7e7b;
            11'd915: table_out = 36'hfb8488746;
            11'd916: table_out = 36'hfb8648df1;
            11'd917: table_out = 36'hfb880927b;
            11'd918: table_out = 36'hfb89c94e5;
            11'd919: table_out = 36'hfb8b8952f;
            11'd920: table_out = 36'hfb8d4935b;
            11'd921: table_out = 36'hfb8f08f67;
            11'd922: table_out = 36'hfb90c8954;
            11'd923: table_out = 36'hfb9288124;
            11'd924: table_out = 36'hfb94476d5;
            11'd925: table_out = 36'hfb9606a68;
            11'd926: table_out = 36'hfb97c5bde;
            11'd927: table_out = 36'hfb9984b37;
            11'd928: table_out = 36'hfb9b43874;
            11'd929: table_out = 36'hfb9d02393;
            11'd930: table_out = 36'hfb9ec0c97;
            11'd931: table_out = 36'hfba07f37f;
            11'd932: table_out = 36'hfba23d84c;
            11'd933: table_out = 36'hfba3fbafd;
            11'd934: table_out = 36'hfba5b9b93;
            11'd935: table_out = 36'hfba777a0f;
            11'd936: table_out = 36'hfba935671;
            11'd937: table_out = 36'hfbaaf30b9;
            11'd938: table_out = 36'hfbacb08e7;
            11'd939: table_out = 36'hfbae6defc;
            11'd940: table_out = 36'hfbb02b2f8;
            11'd941: table_out = 36'hfbb1e84dc;
            11'd942: table_out = 36'hfbb3a54a7;
            11'd943: table_out = 36'hfbb56225a;
            11'd944: table_out = 36'hfbb71edf6;
            11'd945: table_out = 36'hfbb8db77a;
            11'd946: table_out = 36'hfbba97ee7;
            11'd947: table_out = 36'hfbbc5443e;
            11'd948: table_out = 36'hfbbe1077e;
            11'd949: table_out = 36'hfbbfcc8a8;
            11'd950: table_out = 36'hfbc1887bc;
            11'd951: table_out = 36'hfbc3444bb;
            11'd952: table_out = 36'hfbc4fffa4;
            11'd953: table_out = 36'hfbc6bb879;
            11'd954: table_out = 36'hfbc876f39;
            11'd955: table_out = 36'hfbca323e5;
            11'd956: table_out = 36'hfbcbed67d;
            11'd957: table_out = 36'hfbcda8701;
            11'd958: table_out = 36'hfbcf63573;
            11'd959: table_out = 36'hfbd11e1d1;
            11'd960: table_out = 36'hfbd2d8c1c;
            11'd961: table_out = 36'hfbd493455;
            11'd962: table_out = 36'hfbd64da7c;
            11'd963: table_out = 36'hfbd807e92;
            11'd964: table_out = 36'hfbd9c2096;
            11'd965: table_out = 36'hfbdb7c088;
            11'd966: table_out = 36'hfbdd35e6a;
            11'd967: table_out = 36'hfbdeefa3c;
            11'd968: table_out = 36'hfbe0a93fd;
            11'd969: table_out = 36'hfbe262baf;
            11'd970: table_out = 36'hfbe41c151;
            11'd971: table_out = 36'hfbe5d54e3;
            11'd972: table_out = 36'hfbe78e667;
            11'd973: table_out = 36'hfbe9475dc;
            11'd974: table_out = 36'hfbeb00342;
            11'd975: table_out = 36'hfbecb8e9b;
            11'd976: table_out = 36'hfbee717e6;
            11'd977: table_out = 36'hfbf029f23;
            11'd978: table_out = 36'hfbf1e2454;
            11'd979: table_out = 36'hfbf39a777;
            11'd980: table_out = 36'hfbf55288e;
            11'd981: table_out = 36'hfbf70a799;
            11'd982: table_out = 36'hfbf8c2498;
            11'd983: table_out = 36'hfbfa79f8b;
            11'd984: table_out = 36'hfbfc31873;
            11'd985: table_out = 36'hfbfde8f50;
            11'd986: table_out = 36'hfbffa0423;
            11'd987: table_out = 36'hfc01576eb;
            11'd988: table_out = 36'hfc030e7a9;
            11'd989: table_out = 36'hfc04c565d;
            11'd990: table_out = 36'hfc067c308;
            11'd991: table_out = 36'hfc0832da9;
            11'd992: table_out = 36'hfc09e9642;
            11'd993: table_out = 36'hfc0b9fcd2;
            11'd994: table_out = 36'hfc0d5615a;
            11'd995: table_out = 36'hfc0f0c3d9;
            11'd996: table_out = 36'hfc10c2452;
            11'd997: table_out = 36'hfc12782c3;
            11'd998: table_out = 36'hfc142df2c;
            11'd999: table_out = 36'hfc15e398f;
            11'd1000: table_out = 36'hfc17991ec;
            11'd1001: table_out = 36'hfc194e842;
            11'd1002: table_out = 36'hfc1b03c93;
            11'd1003: table_out = 36'hfc1cb8ede;
            11'd1004: table_out = 36'hfc1e6df24;
            11'd1005: table_out = 36'hfc2022d64;
            11'd1006: table_out = 36'hfc21d79a1;
            11'd1007: table_out = 36'hfc238c3d8;
            11'd1008: table_out = 36'hfc2540c0c;
            11'd1009: table_out = 36'hfc26f523c;
            11'd1010: table_out = 36'hfc28a9668;
            11'd1011: table_out = 36'hfc2a5d892;
            11'd1012: table_out = 36'hfc2c118b8;
            11'd1013: table_out = 36'hfc2dc56dc;
            11'd1014: table_out = 36'hfc2f792fe;
            11'd1015: table_out = 36'hfc312cd1d;
            11'd1016: table_out = 36'hfc32e053b;
            11'd1017: table_out = 36'hfc3493b57;
            11'd1018: table_out = 36'hfc3646f73;
            11'd1019: table_out = 36'hfc37fa18d;
            11'd1020: table_out = 36'hfc39ad1a8;
            11'd1021: table_out = 36'hfc3b5ffc1;
            11'd1022: table_out = 36'hfc3d12bdb;
            11'd1023: table_out = 36'hfc3ec55f6;
            11'd1024: table_out = 36'hfc4077e11;
            11'd1025: table_out = 36'hfc422a42d;
            11'd1026: table_out = 36'hfc43dc84a;
            11'd1027: table_out = 36'hfc458ea68;
            11'd1028: table_out = 36'hfc4740a89;
            11'd1029: table_out = 36'hfc48f28ac;
            11'd1030: table_out = 36'hfc4aa44d1;
            11'd1031: table_out = 36'hfc4c55ef9;
            11'd1032: table_out = 36'hfc4e07724;
            11'd1033: table_out = 36'hfc4fb8d52;
            11'd1034: table_out = 36'hfc516a184;
            11'd1035: table_out = 36'hfc531b3b9;
            11'd1036: table_out = 36'hfc54cc3f3;
            11'd1037: table_out = 36'hfc567d231;
            11'd1038: table_out = 36'hfc582de74;
            11'd1039: table_out = 36'hfc59de8bd;
            11'd1040: table_out = 36'hfc5b8f10a;
            11'd1041: table_out = 36'hfc5d3f75d;
            11'd1042: table_out = 36'hfc5eefbb6;
            11'd1043: table_out = 36'hfc609fe15;
            11'd1044: table_out = 36'hfc624fe7b;
            11'd1045: table_out = 36'hfc63ffce7;
            11'd1046: table_out = 36'hfc65af95b;
            11'd1047: table_out = 36'hfc675f3d6;
            11'd1048: table_out = 36'hfc690ec58;
            11'd1049: table_out = 36'hfc6abe2e3;
            11'd1050: table_out = 36'hfc6c6d775;
            11'd1051: table_out = 36'hfc6e1ca11;
            11'd1052: table_out = 36'hfc6fcbab5;
            11'd1053: table_out = 36'hfc717a962;
            11'd1054: table_out = 36'hfc7329618;
            11'd1055: table_out = 36'hfc74d80d8;
            11'd1056: table_out = 36'hfc76869a2;
            11'd1057: table_out = 36'hfc7835076;
            11'd1058: table_out = 36'hfc79e3555;
            11'd1059: table_out = 36'hfc7b9183f;
            11'd1060: table_out = 36'hfc7d3f933;
            11'd1061: table_out = 36'hfc7eed833;
            11'd1062: table_out = 36'hfc809b53f;
            11'd1063: table_out = 36'hfc8249057;
            11'd1064: table_out = 36'hfc83f697b;
            11'd1065: table_out = 36'hfc85a40ab;
            11'd1066: table_out = 36'hfc87515e8;
            11'd1067: table_out = 36'hfc88fe932;
            11'd1068: table_out = 36'hfc8aaba8a;
            11'd1069: table_out = 36'hfc8c589ef;
            11'd1070: table_out = 36'hfc8e05762;
            11'd1071: table_out = 36'hfc8fb22e3;
            11'd1072: table_out = 36'hfc915ec73;
            11'd1073: table_out = 36'hfc930b412;
            11'd1074: table_out = 36'hfc94b79bf;
            11'd1075: table_out = 36'hfc9663d7c;
            11'd1076: table_out = 36'hfc980ff49;
            11'd1077: table_out = 36'hfc99bbf25;
            11'd1078: table_out = 36'hfc9b67d12;
            11'd1079: table_out = 36'hfc9d1390f;
            11'd1080: table_out = 36'hfc9ebf31c;
            11'd1081: table_out = 36'hfca06ab3b;
            11'd1082: table_out = 36'hfca21616b;
            11'd1083: table_out = 36'hfca3c15ad;
            11'd1084: table_out = 36'hfca56c800;
            11'd1085: table_out = 36'hfca717866;
            11'd1086: table_out = 36'hfca8c26de;
            11'd1087: table_out = 36'hfcaa6d369;
            11'd1088: table_out = 36'hfcac17e06;
            11'd1089: table_out = 36'hfcadc26b7;
            11'd1090: table_out = 36'hfcaf6cd7c;
            11'd1091: table_out = 36'hfcb117254;
            11'd1092: table_out = 36'hfcb2c1540;
            11'd1093: table_out = 36'hfcb46b641;
            11'd1094: table_out = 36'hfcb615556;
            11'd1095: table_out = 36'hfcb7bf280;
            11'd1096: table_out = 36'hfcb968dc0;
            11'd1097: table_out = 36'hfcbb12715;
            11'd1098: table_out = 36'hfcbcbbe7f;
            11'd1099: table_out = 36'hfcbe65400;
            11'd1100: table_out = 36'hfcc00e796;
            11'd1101: table_out = 36'hfcc1b7944;
            11'd1102: table_out = 36'hfcc360908;
            11'd1103: table_out = 36'hfcc5096e4;
            11'd1104: table_out = 36'hfcc6b22d6;
            11'd1105: table_out = 36'hfcc85ace1;
            11'd1106: table_out = 36'hfcca03503;
            11'd1107: table_out = 36'hfccbabb3e;
            11'd1108: table_out = 36'hfccd53f91;
            11'd1109: table_out = 36'hfccefc1fc;
            11'd1110: table_out = 36'hfcd0a4281;
            11'd1111: table_out = 36'hfcd24c11f;
            11'd1112: table_out = 36'hfcd3f3dd7;
            11'd1113: table_out = 36'hfcd59b8a8;
            11'd1114: table_out = 36'hfcd743194;
            11'd1115: table_out = 36'hfcd8ea89a;
            11'd1116: table_out = 36'hfcda91dbb;
            11'd1117: table_out = 36'hfcdc390f6;
            11'd1118: table_out = 36'hfcdde024d;
            11'd1119: table_out = 36'hfcdf871bf;
            11'd1120: table_out = 36'hfce12df4d;
            11'd1121: table_out = 36'hfce2d4af7;
            11'd1122: table_out = 36'hfce47b4be;
            11'd1123: table_out = 36'hfce621ca1;
            11'd1124: table_out = 36'hfce7c82a0;
            11'd1125: table_out = 36'hfce96e6bd;
            11'd1126: table_out = 36'hfceb148f7;
            11'd1127: table_out = 36'hfcecba94f;
            11'd1128: table_out = 36'hfcee607c5;
            11'd1129: table_out = 36'hfcf006459;
            11'd1130: table_out = 36'hfcf1abf0b;
            11'd1131: table_out = 36'hfcf3517dc;
            11'd1132: table_out = 36'hfcf4f6ecc;
            11'd1133: table_out = 36'hfcf69c3dc;
            11'd1134: table_out = 36'hfcf84170a;
            11'd1135: table_out = 36'hfcf9e6859;
            11'd1136: table_out = 36'hfcfb8b7c8;
            11'd1137: table_out = 36'hfcfd30556;
            11'd1138: table_out = 36'hfcfed5106;
            11'd1139: table_out = 36'hfd0079ad6;
            11'd1140: table_out = 36'hfd021e2c8;
            11'd1141: table_out = 36'hfd03c28db;
            11'd1142: table_out = 36'hfd0566d0f;
            11'd1143: table_out = 36'hfd070af66;
            11'd1144: table_out = 36'hfd08aefde;
            11'd1145: table_out = 36'hfd0a52e79;
            11'd1146: table_out = 36'hfd0bf6b37;
            11'd1147: table_out = 36'hfd0d9a618;
            11'd1148: table_out = 36'hfd0f3df1c;
            11'd1149: table_out = 36'hfd10e1643;
            11'd1150: table_out = 36'hfd1284b8e;
            11'd1151: table_out = 36'hfd1427efe;
            11'd1152: table_out = 36'hfd15cb091;
            11'd1153: table_out = 36'hfd176e049;
            11'd1154: table_out = 36'hfd1910e26;
            11'd1155: table_out = 36'hfd1ab3a28;
            11'd1156: table_out = 36'hfd1c56450;
            11'd1157: table_out = 36'hfd1df8c9d;
            11'd1158: table_out = 36'hfd1f9b30f;
            11'd1159: table_out = 36'hfd213d7a8;
            11'd1160: table_out = 36'hfd22dfa68;
            11'd1161: table_out = 36'hfd2481b4e;
            11'd1162: table_out = 36'hfd2623a5b;
            11'd1163: table_out = 36'hfd27c578f;
            11'd1164: table_out = 36'hfd29672ea;
            11'd1165: table_out = 36'hfd2b08c6e;
            11'd1166: table_out = 36'hfd2caa419;
            11'd1167: table_out = 36'hfd2e4b9ec;
            11'd1168: table_out = 36'hfd2fecde8;
            11'd1169: table_out = 36'hfd318e00d;
            11'd1170: table_out = 36'hfd332f05b;
            11'd1171: table_out = 36'hfd34cfed2;
            11'd1172: table_out = 36'hfd3670b72;
            11'd1173: table_out = 36'hfd381163d;
            11'd1174: table_out = 36'hfd39b1f31;
            11'd1175: table_out = 36'hfd3b52650;
            11'd1176: table_out = 36'hfd3cf2b99;
            11'd1177: table_out = 36'hfd3e92f0d;
            11'd1178: table_out = 36'hfd40330ac;
            11'd1179: table_out = 36'hfd41d3076;
            11'd1180: table_out = 36'hfd4372e6c;
            11'd1181: table_out = 36'hfd4512a8e;
            11'd1182: table_out = 36'hfd46b24dc;
            11'd1183: table_out = 36'hfd4851d56;
            11'd1184: table_out = 36'hfd49f13fd;
            11'd1185: table_out = 36'hfd4b908d1;
            11'd1186: table_out = 36'hfd4d2fbd2;
            11'd1187: table_out = 36'hfd4eced00;
            11'd1188: table_out = 36'hfd506dc5c;
            11'd1189: table_out = 36'hfd520c9e6;
            11'd1190: table_out = 36'hfd53ab59e;
            11'd1191: table_out = 36'hfd5549f85;
            11'd1192: table_out = 36'hfd56e879a;
            11'd1193: table_out = 36'hfd5886dde;
            11'd1194: table_out = 36'hfd5a25251;
            11'd1195: table_out = 36'hfd5bc34f4;
            11'd1196: table_out = 36'hfd5d615c6;
            11'd1197: table_out = 36'hfd5eff4c8;
            11'd1198: table_out = 36'hfd609d1fb;
            11'd1199: table_out = 36'hfd623ad5d;
            11'd1200: table_out = 36'hfd63d86f1;
            11'd1201: table_out = 36'hfd6575eb6;
            11'd1202: table_out = 36'hfd67134ab;
            11'd1203: table_out = 36'hfd68b08d3;
            11'd1204: table_out = 36'hfd6a4db2c;
            11'd1205: table_out = 36'hfd6beabb6;
            11'd1206: table_out = 36'hfd6d87a74;
            11'd1207: table_out = 36'hfd6f24763;
            11'd1208: table_out = 36'hfd70c1285;
            11'd1209: table_out = 36'hfd725dbdb;
            11'd1210: table_out = 36'hfd73fa363;
            11'd1211: table_out = 36'hfd759691f;
            11'd1212: table_out = 36'hfd7732d0f;
            11'd1213: table_out = 36'hfd78cef32;
            11'd1214: table_out = 36'hfd7a6af8a;
            11'd1215: table_out = 36'hfd7c06e17;
            11'd1216: table_out = 36'hfd7da2ad8;
            11'd1217: table_out = 36'hfd7f3e5ce;
            11'd1218: table_out = 36'hfd80d9ef9;
            11'd1219: table_out = 36'hfd827565a;
            11'd1220: table_out = 36'hfd8410bf1;
            11'd1221: table_out = 36'hfd85abfbd;
            11'd1222: table_out = 36'hfd87471c0;
            11'd1223: table_out = 36'hfd88e21f9;
            11'd1224: table_out = 36'hfd8a7d069;
            11'd1225: table_out = 36'hfd8c17d10;
            11'd1226: table_out = 36'hfd8db27ee;
            11'd1227: table_out = 36'hfd8f4d103;
            11'd1228: table_out = 36'hfd90c10bb;
            default: table_out = 36'b0;
        endcase
    end

endmodule