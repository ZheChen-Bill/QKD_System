
//226 * 36
//36 word length
//32 fraction length

module ln_lam_1_lam_table(
    input [8-1:0] index, //0~255
    output reg [36-1:0] table_out //36 word length, 32 fraction length
);


    always@(*) begin
        case(index)
            8'd0: table_out = 36'hd1f706e0b;
            8'd1: table_out = 36'hd1e75b0cc;
            8'd2: table_out = 36'hd1d79d938;
            8'd3: table_out = 36'hd1c7ce4fe;
            8'd4: table_out = 36'hd1b7ed1c5;
            8'd5: table_out = 36'hd1a7f9d2e;
            8'd6: table_out = 36'hd197f44d2;
            8'd7: table_out = 36'hd187dc641;
            8'd8: table_out = 36'hd177b1f05;
            8'd9: table_out = 36'hd16774c9e;
            8'd10: table_out = 36'hd15724c85;
            8'd11: table_out = 36'hd146c1c2b;
            8'd12: table_out = 36'hd1364b8f9;
            8'd13: table_out = 36'hd125c204d;
            8'd14: table_out = 36'hd11524f7f;
            8'd15: table_out = 36'hd104743dd;
            8'd16: table_out = 36'hd0f3afaac;
            8'd17: table_out = 36'hd0e2d7127;
            8'd18: table_out = 36'hd0d1ea482;
            8'd19: table_out = 36'hd0c0e91e5;
            8'd20: table_out = 36'hd0afd3671;
            8'd21: table_out = 36'hd09ea8f3a;
            8'd22: table_out = 36'hd08d6994c;
            8'd23: table_out = 36'hd07c151a8;
            8'd24: table_out = 36'hd06aab546;
            8'd25: table_out = 36'hd0592c112;
            8'd26: table_out = 36'hd047971ee;
            8'd27: table_out = 36'hd035ec4b0;
            8'd28: table_out = 36'hd0242b624;
            8'd29: table_out = 36'hd0125430a;
            8'd30: table_out = 36'hd00066818;
            8'd31: table_out = 36'hcfee621f5;
            8'd32: table_out = 36'hcfdc46d3f;
            8'd33: table_out = 36'hcfca14687;
            8'd34: table_out = 36'hcfb7caa50;
            8'd35: table_out = 36'hcfa569512;
            8'd36: table_out = 36'hcf92f0338;
            8'd37: table_out = 36'hcf805f11f;
            8'd38: table_out = 36'hcf6db5b18;
            8'd39: table_out = 36'hcf5af3d64;
            8'd40: table_out = 36'hcf4819437;
            8'd41: table_out = 36'hcf3525bb8;
            8'd42: table_out = 36'hcf2218ffe;
            8'd43: table_out = 36'hcf0ef2d12;
            8'd44: table_out = 36'hcefbb2eed;
            8'd45: table_out = 36'hcee85917b;
            8'd46: table_out = 36'hced4e5094;
            8'd47: table_out = 36'hcec156804;
            8'd48: table_out = 36'hceadad385;
            8'd49: table_out = 36'hce99e8ec1;
            8'd50: table_out = 36'hce860954f;
            8'd51: table_out = 36'hce720e2b7;
            8'd52: table_out = 36'hce5df726e;
            8'd53: table_out = 36'hce49c3fd8;
            8'd54: table_out = 36'hce3574644;
            8'd55: table_out = 36'hce21080f2;
            8'd56: table_out = 36'hce0c7eb0c;
            8'd57: table_out = 36'hcdf7d7fa8;
            8'd58: table_out = 36'hcde3139ca;
            8'd59: table_out = 36'hcdce3145f;
            8'd60: table_out = 36'hcdb930a42;
            8'd61: table_out = 36'hcda411636;
            8'd62: table_out = 36'hcd8ed32ea;
            8'd63: table_out = 36'hcd7975af5;
            8'd64: table_out = 36'hcd63f88d8;
            8'd65: table_out = 36'hcd4e5b6fd;
            8'd66: table_out = 36'hcd389dfb5;
            8'd67: table_out = 36'hcd22bfd3a;
            8'd68: table_out = 36'hcd0cc09ab;
            8'd69: table_out = 36'hccf69ff10;
            8'd70: table_out = 36'hcce05d756;
            8'd71: table_out = 36'hccc9f8c4e;
            8'd72: table_out = 36'hccb3717af;
            8'd73: table_out = 36'hcc9cc7313;
            8'd74: table_out = 36'hcc85f97fa;
            8'd75: table_out = 36'hcc6f07fc3;
            8'd76: table_out = 36'hcc57f23b1;
            8'd77: table_out = 36'hcc40b7cea;
            8'd78: table_out = 36'hcc2958471;
            8'd79: table_out = 36'hcc11d332b;
            8'd80: table_out = 36'hcbfa281dc;
            8'd81: table_out = 36'hcbe256926;
            8'd82: table_out = 36'hcbca5e188;
            8'd83: table_out = 36'hcbb23e35f;
            8'd84: table_out = 36'hcb99f66e1;
            8'd85: table_out = 36'hcb8186423;
            8'd86: table_out = 36'hcb68ed310;
            8'd87: table_out = 36'hcb502ab6d;
            8'd88: table_out = 36'hcb373e4d8;
            8'd89: table_out = 36'hcb1e276c5;
            8'd90: table_out = 36'hcb04e587f;
            8'd91: table_out = 36'hcaeb78123;
            8'd92: table_out = 36'hcad1de7a5;
            8'd93: table_out = 36'hcab8182ca;
            8'd94: table_out = 36'hca9e24927;
            8'd95: table_out = 36'hca8403124;
            8'd96: table_out = 36'hca69b30f5;
            8'd97: table_out = 36'hca4f33e9d;
            8'd98: table_out = 36'hca3484fea;
            8'd99: table_out = 36'hca19a5a76;
            8'd100: table_out = 36'hc9fe953a3;
            8'd101: table_out = 36'hc9e35309b;
            8'd102: table_out = 36'hc9c7de64f;
            8'd103: table_out = 36'hc9ac36973;
            8'd104: table_out = 36'hc9905ae7f;
            8'd105: table_out = 36'hc9744a9ab;
            8'd106: table_out = 36'hc95804eef;
            8'd107: table_out = 36'hc93b89200;
            8'd108: table_out = 36'hc91ed6650;
            8'd109: table_out = 36'hc901ebf08;
            8'd110: table_out = 36'hc8e4c8f0a;
            8'd111: table_out = 36'hc8c76c8ed;
            8'd112: table_out = 36'hc8a9d5efb;
            8'd113: table_out = 36'hc88c0432d;
            8'd114: table_out = 36'hc86df672e;
            8'd115: table_out = 36'hc84fabc50;
            8'd116: table_out = 36'hc83123393;
            8'd117: table_out = 36'hc8125bd9a;
            8'd118: table_out = 36'hc7f354aad;
            8'd119: table_out = 36'hc7d40cab5;
            8'd120: table_out = 36'hc7b482d38;
            8'd121: table_out = 36'hc794b6156;
            8'd122: table_out = 36'hc774a55c8;
            8'd123: table_out = 36'hc7544f8db;
            8'd124: table_out = 36'hc733b3869;
            8'd125: table_out = 36'hc712d01dd;
            8'd126: table_out = 36'hc6f1a4229;
            8'd127: table_out = 36'hc6d02e5c2;
            8'd128: table_out = 36'hc6ae6d8a0;
            8'd129: table_out = 36'hc68c60636;
            8'd130: table_out = 36'hc66a0596f;
            8'd131: table_out = 36'hc6475bcaa;
            8'd132: table_out = 36'hc624619b2;
            8'd133: table_out = 36'hc601159bb;
            8'd134: table_out = 36'hc5dd7655e;
            8'd135: table_out = 36'hc5b982490;
            8'd136: table_out = 36'hc59537e9f;
            8'd137: table_out = 36'hc57095a29;
            8'd138: table_out = 36'hc54b99d19;
            8'd139: table_out = 36'hc52642c9e;
            8'd140: table_out = 36'hc5008ed22;
            8'd141: table_out = 36'hc4da7c248;
            8'd142: table_out = 36'hc4b408edf;
            8'd143: table_out = 36'hc48d334dd;
            8'd144: table_out = 36'hc465f9553;
            8'd145: table_out = 36'hc43e59069;
            8'd146: table_out = 36'hc41650550;
            8'd147: table_out = 36'hc3eddd23c;
            8'd148: table_out = 36'hc3c4fd454;
            8'd149: table_out = 36'hc39bae7ad;
            8'd150: table_out = 36'hc371ee73c;
            8'd151: table_out = 36'hc347bacc9;
            8'd152: table_out = 36'hc31d110e2;
            8'd153: table_out = 36'hc2f1eeacf;
            8'd154: table_out = 36'hc2c651085;
            8'd155: table_out = 36'hc29a35693;
            8'd156: table_out = 36'hc26d99015;
            8'd157: table_out = 36'hc24078ea3;
            8'd158: table_out = 36'hc212d223d;
            8'd159: table_out = 36'hc1e4a193d;
            8'd160: table_out = 36'hc1b5e403e;
            8'd161: table_out = 36'hc1869620a;
            8'd162: table_out = 36'hc156b4784;
            8'd163: table_out = 36'hc1263b78e;
            8'd164: table_out = 36'hc0f5276f1;
            8'd165: table_out = 36'hc0c374846;
            8'd166: table_out = 36'hc0911ebd3;
            8'd167: table_out = 36'hc05e21f74;
            8'd168: table_out = 36'hc02a79e73;
            8'd169: table_out = 36'hbff622170;
            8'd170: table_out = 36'hbfc115e33;
            8'd171: table_out = 36'hbf8b5078c;
            8'd172: table_out = 36'hbf54ccd26;
            8'd173: table_out = 36'hbf1d85b5c;
            8'd174: table_out = 36'hbee575b0b;
            8'd175: table_out = 36'hbeac9715c;
            8'd176: table_out = 36'hbe72e3f91;
            8'd177: table_out = 36'hbe38562ca;
            8'd178: table_out = 36'hbdfce73c7;
            8'd179: table_out = 36'hbdc0906a1;
            8'd180: table_out = 36'hbd834aa87;
            8'd181: table_out = 36'hbd450e96e;
            8'd182: table_out = 36'hbd05d47bb;
            8'd183: table_out = 36'hbcc5943ed;
            8'd184: table_out = 36'hbc8445637;
            8'd185: table_out = 36'hbc41df015;
            8'd186: table_out = 36'hbbfe57be0;
            8'd187: table_out = 36'hbbb9a5c47;
            8'd188: table_out = 36'hbb73bebd2;
            8'd189: table_out = 36'hbb2c97c46;
            8'd190: table_out = 36'hbae42560a;
            8'd191: table_out = 36'hba9a5b774;
            8'd192: table_out = 36'hba4f2d40d;
            8'd193: table_out = 36'hba028d3ba;
            8'd194: table_out = 36'hb9b46d1da;
            8'd195: table_out = 36'hb964bdc4b;
            8'd196: table_out = 36'hb9136f24b;
            8'd197: table_out = 36'hb8c070351;
            8'd198: table_out = 36'hb86baedb0;
            8'd199: table_out = 36'hb81517d26;
            8'd200: table_out = 36'hb7bc96938;
            8'd201: table_out = 36'hb76215369;
            8'd202: table_out = 36'hb7057c52e;
            8'd203: table_out = 36'hb6a6b2db7;
            8'd204: table_out = 36'hb6459df63;
            8'd205: table_out = 36'hb5e220cf0;
            8'd206: table_out = 36'hb57c1c64c;
            8'd207: table_out = 36'hb5136f4fa;
            8'd208: table_out = 36'hb4a7f5803;
            8'd209: table_out = 36'hb43987f52;
            8'd210: table_out = 36'hb3c7fc673;
            8'd211: table_out = 36'hb35324e87;
            8'd212: table_out = 36'hb2dacf75a;
            8'd213: table_out = 36'hb25ec5765;
            8'd214: table_out = 36'hb1decb290;
            8'd215: table_out = 36'hb15a9ef76;
            8'd216: table_out = 36'hb0d1f8ad5;
            8'd217: table_out = 36'hb044888d3;
            8'd218: table_out = 36'hafb1f6398;
            8'd219: table_out = 36'haf19df6a9;
            8'd220: table_out = 36'hae7bd663e;
            8'd221: table_out = 36'hadd76019d;
            8'd222: table_out = 36'had2bf1f31;
            8'd223: table_out = 36'hac78ef0c3;
            8'd224: table_out = 36'habbda4d95;
            8'd225: table_out = 36'hab4150edf;
            default: table_out = 36'b0;
        endcase
    end

endmodule